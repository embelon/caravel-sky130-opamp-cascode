* NGSPICE file created from top_ew_algofoogle.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

.subckt top_ew_algofoogle i_clk i_debug_map_overlay i_debug_trace_overlay i_debug_vec_overlay
+ i_gpout0_sel[0] i_gpout0_sel[1] i_gpout0_sel[2] i_gpout0_sel[3] i_gpout0_sel[4]
+ i_gpout0_sel[5] i_gpout1_sel[0] i_gpout1_sel[1] i_gpout1_sel[2] i_gpout1_sel[3]
+ i_gpout1_sel[4] i_gpout1_sel[5] i_gpout2_sel[0] i_gpout2_sel[1] i_gpout2_sel[2]
+ i_gpout2_sel[3] i_gpout2_sel[4] i_gpout2_sel[5] i_gpout3_sel[0] i_gpout3_sel[1]
+ i_gpout3_sel[2] i_gpout3_sel[3] i_gpout3_sel[4] i_gpout3_sel[5] i_gpout4_sel[0]
+ i_gpout4_sel[1] i_gpout4_sel[2] i_gpout4_sel[3] i_gpout4_sel[4] i_gpout4_sel[5]
+ i_gpout5_sel[0] i_gpout5_sel[1] i_gpout5_sel[2] i_gpout5_sel[3] i_gpout5_sel[4]
+ i_gpout5_sel[5] i_la_invalid i_mode[0] i_mode[1] i_mode[2] i_reg_csb i_reg_mosi
+ i_reg_sclk i_reset_lock_a i_reset_lock_b i_tex_in[0] i_tex_in[1] i_tex_in[2] i_tex_in[3]
+ i_vec_csb i_vec_mosi i_vec_sclk o_gpout[0] o_gpout[1] o_gpout[2] o_gpout[3] o_gpout[4]
+ o_gpout[5] o_hsync o_reset o_rgb[0] o_rgb[10] o_rgb[11] o_rgb[12] o_rgb[13] o_rgb[14]
+ o_rgb[15] o_rgb[16] o_rgb[17] o_rgb[18] o_rgb[19] o_rgb[1] o_rgb[20] o_rgb[21] o_rgb[22]
+ o_rgb[23] o_rgb[2] o_rgb[3] o_rgb[4] o_rgb[5] o_rgb[6] o_rgb[7] o_rgb[8] o_rgb[9]
+ o_tex_csb o_tex_oeb0 o_tex_out0 o_tex_sclk o_vsync ones[0] ones[10] ones[11] ones[12]
+ ones[13] ones[14] ones[15] ones[1] ones[2] ones[3] ones[4] ones[5] ones[6] ones[7]
+ ones[8] ones[9] vccd1 vssd1 zeros[0] zeros[10] zeros[11] zeros[12] zeros[13] zeros[14]
+ zeros[15] zeros[1] zeros[2] zeros[3] zeros[4] zeros[5] zeros[6] zeros[7] zeros[8]
+ zeros[9]
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18869_ rbzero.wall_tracer.trackDistY\[9\] _02542_ _02398_ vssd1 vssd1 vccd1 vccd1
+ _02543_ sky130_fd_sc_hd__mux2_1
XFILLER_28_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20900_ clknet_leaf_85_i_clk _00669_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_20831_ clknet_leaf_51_i_clk _00600_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20762_ clknet_leaf_46_i_clk _00531_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_195_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20693_ clknet_leaf_58_i_clk _00477_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21314_ net235 _01083_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_164_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21245_ clknet_leaf_91_i_clk _01014_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_104_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21176_ clknet_leaf_5_i_clk _00945_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20127_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__buf_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11900_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _04290_ vssd1 vssd1 vccd1 vccd1 _04676_
+ sky130_fd_sc_hd__mux2_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12880_ rbzero.wall_tracer.visualWallDist\[-1\] _05571_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05617_ sky130_fd_sc_hd__a21o_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _04605_ _04606_ _04607_ _04266_ _04229_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__o221a_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14550_ _07259_ _07266_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__xnor2_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _04129_ vssd1 vssd1 vccd1 vccd1 _04540_
+ sky130_fd_sc_hd__mux2_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ _06201_ _06204_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__or2_1
XFILLER_198_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10713_ rbzero.tex_g1\[1\] rbzero.tex_g1\[2\] _03691_ vssd1 vssd1 vccd1 vccd1 _03698_
+ sky130_fd_sc_hd__mux2_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _07216_ _07217_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__nor2_2
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11693_ rbzero.debug_overlay.vplaneY\[-4\] _04464_ _04460_ rbzero.debug_overlay.vplaneY\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a22o_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16220_ _08860_ _08864_ vssd1 vssd1 vccd1 vccd1 _08865_ sky130_fd_sc_hd__or2_1
X_13432_ _06156_ _06167_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__and2_1
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10644_ rbzero.tex_g1\[34\] rbzero.tex_g1\[35\] _03658_ vssd1 vssd1 vccd1 vccd1 _03662_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _08795_ _08792_ vssd1 vssd1 vccd1 vccd1 _08796_ sky130_fd_sc_hd__xnor2_1
X_10575_ _03625_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13363_ _05823_ _05973_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__or2_1
XFILLER_166_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15102_ _07757_ _07758_ _07759_ _07760_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__nand4_2
X_12314_ net27 vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__clkbuf_4
XFILLER_177_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16082_ _08283_ _08491_ vssd1 vssd1 vccd1 vccd1 _08727_ sky130_fd_sc_hd__or2_1
XFILLER_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13294_ _05975_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__clkbuf_4
XFILLER_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15033_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__nor2_1
X_19910_ rbzero.pov.ready_buffer\[50\] _03141_ _03192_ _03210_ vssd1 vssd1 vccd1 vccd1
+ _03211_ sky130_fd_sc_hd__a211o_1
X_12245_ net41 _04962_ _04978_ net43 net17 vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__a221o_1
XFILLER_142_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12176_ _04907_ net10 _04944_ _04946_ net11 vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__a311o_1
X_19841_ rbzero.pov.ready_buffer\[64\] _07948_ _03146_ vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11127_ rbzero.wall_tracer.visualWallDist\[8\] rbzero.wall_tracer.visualWallDist\[7\]
+ rbzero.wall_tracer.visualWallDist\[6\] rbzero.wall_tracer.visualWallDist\[5\] vssd1
+ vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__or4_1
X_16984_ _09620_ _09623_ vssd1 vssd1 vccd1 vccd1 _09624_ sky130_fd_sc_hd__nand2_1
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19772_ rbzero.pov.spi_buffer\[59\] rbzero.pov.spi_buffer\[60\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03115_ sky130_fd_sc_hd__mux2_1
XFILLER_110_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15935_ _08129_ _08579_ vssd1 vssd1 vccd1 vccd1 _08580_ sky130_fd_sc_hd__or2_2
XFILLER_77_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18723_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.stepDistY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__nand2_1
X_11058_ rbzero.tex_b0\[30\] rbzero.tex_b0\[29\] _03876_ vssd1 vssd1 vccd1 vccd1 _03879_
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18654_ _02330_ _02349_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__xnor2_1
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ _08510_ _08466_ vssd1 vssd1 vccd1 vccd1 _08511_ sky130_fd_sc_hd__xnor2_4
XFILLER_149_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17605_ _10167_ _10170_ vssd1 vssd1 vccd1 vccd1 _10171_ sky130_fd_sc_hd__xnor2_2
X_14817_ _07487_ _07456_ _07544_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__a21o_1
X_18585_ _02269_ _02270_ _02281_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a21oi_1
Xtop_ew_algofoogle_120 vssd1 vssd1 vccd1 vccd1 ones[14] top_ew_algofoogle_120/LO sky130_fd_sc_hd__conb_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15797_ _08382_ _08388_ vssd1 vssd1 vccd1 vccd1 _08442_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17536_ _09126_ _09674_ vssd1 vssd1 vccd1 vccd1 _10102_ sky130_fd_sc_hd__nor2_1
XFILLER_33_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14748_ _05814_ _07472_ _07482_ _07459_ vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__o211a_1
XFILLER_205_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17467_ _10030_ _10031_ _10029_ _09902_ vssd1 vssd1 vccd1 vccd1 _10034_ sky130_fd_sc_hd__o211a_1
X_14679_ _07343_ _07344_ _07346_ _07378_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__o211a_1
XFILLER_149_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20140__170 clknet_1_0__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__inv_2
X_19206_ _02750_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__clkbuf_1
X_16418_ rbzero.debug_overlay.playerY\[-6\] rbzero.debug_overlay.playerX\[-6\] _07895_
+ vssd1 vssd1 vccd1 vccd1 _09063_ sky130_fd_sc_hd__mux2_1
XFILLER_193_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17398_ _09670_ _09964_ vssd1 vssd1 vccd1 vccd1 _09965_ sky130_fd_sc_hd__xnor2_2
XFILLER_192_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19137_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1
+ _02704_ sky130_fd_sc_hd__and3_1
XFILLER_118_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16349_ _08991_ _08993_ vssd1 vssd1 vccd1 vccd1 _08994_ sky130_fd_sc_hd__xnor2_2
XFILLER_145_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19068_ _02666_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18019_ _10094_ _08423_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__nor2_1
XFILLER_160_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21030_ clknet_leaf_13_i_clk _00799_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20223__245 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__inv_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20814_ clknet_leaf_54_i_clk _00583_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12189__389 _04959_ vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__inv_2
X_20745_ clknet_leaf_44_i_clk _00514_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20676_ clknet_leaf_48_i_clk _00460_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[5\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_7_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03292_ clknet_0__03292_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03292_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10360_ _03510_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12030_ _04140_ _04754_ _04771_ _04787_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__o32a_1
X_21228_ clknet_leaf_17_i_clk _00997_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21159_ clknet_leaf_85_i_clk _00928_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13981_ _06716_ _06717_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__nand2_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15720_ _08363_ _08364_ vssd1 vssd1 vccd1 vccd1 _08365_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_52_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12932_ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__inv_2
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _08288_ _08295_ vssd1 vssd1 vccd1 vccd1 _08296_ sky130_fd_sc_hd__xnor2_4
XFILLER_74_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _05584_ _05586_ _05587_ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__or4b_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _07149_ _07324_ _06176_ _07116_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _01462_ _09703_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__nand2_1
X_11814_ rbzero.color_sky\[2\] rbzero.color_floor\[2\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04592_ sky130_fd_sc_hd__mux2_2
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15582_ _05207_ _08226_ vssd1 vssd1 vccd1 vccd1 _08227_ sky130_fd_sc_hd__nor2_4
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _05534_ _05536_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__or2_1
XFILLER_96_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20198__222 clknet_1_0__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__inv_2
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09890_ sky130_fd_sc_hd__nor2_1
XFILLER_159_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14533_ _07258_ _07050_ _07052_ _07269_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__o31ai_2
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ rbzero.tex_g0\[14\] _04356_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__and2_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17252_ rbzero.wall_tracer.trackDistX\[-10\] _09828_ _05414_ vssd1 vssd1 vccd1 vccd1
+ _09829_ sky130_fd_sc_hd__mux2_1
XFILLER_175_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14464_ _07151_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__inv_2
XFILLER_202_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11676_ _04428_ _04447_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__and2_2
XFILLER_105_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16203_ _08799_ _08798_ vssd1 vssd1 vccd1 vccd1 _08848_ sky130_fd_sc_hd__and2b_1
X_13415_ _06051_ _06090_ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__a21oi_1
X_10627_ rbzero.tex_g1\[42\] rbzero.tex_g1\[43\] _03647_ vssd1 vssd1 vccd1 vccd1 _03653_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17183_ rbzero.traced_texa\[10\] _09770_ _09771_ rbzero.wall_tracer.visualWallDist\[10\]
+ vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__a22o_1
XFILLER_31_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14395_ _07130_ _07131_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__nand2_1
XFILLER_10_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16134_ _08741_ _08753_ vssd1 vssd1 vccd1 vccd1 _08779_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13346_ _06061_ _06067_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__or2_1
X_10558_ _03616_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16065_ _08701_ _08708_ vssd1 vssd1 vccd1 vccd1 _08710_ sky130_fd_sc_hd__nor2_1
X_13277_ _05986_ _06013_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__xnor2_2
X_10489_ _03557_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15016_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.wall_tracer.rayAddendX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__nand2_1
X_12228_ net50 _04978_ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a21oi_1
XFILLER_155_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19824_ _02728_ _02820_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__nor2_1
X_12159_ net11 net10 _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__and3b_1
XFILLER_69_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19755_ rbzero.pov.spi_buffer\[51\] rbzero.pov.spi_buffer\[52\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03106_ sky130_fd_sc_hd__mux2_1
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16967_ _09516_ _09477_ vssd1 vssd1 vccd1 vccd1 _09607_ sky130_fd_sc_hd__or2b_1
X_18706_ _02400_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__clkbuf_1
X_15918_ _08558_ _08562_ vssd1 vssd1 vccd1 vccd1 _08563_ sky130_fd_sc_hd__or2b_1
XFILLER_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16898_ _09410_ _09412_ _09270_ _09409_ vssd1 vssd1 vccd1 vccd1 _09539_ sky130_fd_sc_hd__a2bb2o_1
X_19686_ _03069_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18637_ _02275_ _02276_ _02332_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a21oi_1
X_15849_ _08047_ _08135_ _08491_ _08493_ vssd1 vssd1 vccd1 vccd1 _08494_ sky130_fd_sc_hd__o22ai_4
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18568_ _02263_ _02264_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17519_ _10051_ _10052_ _10084_ vssd1 vssd1 vccd1 vccd1 _10085_ sky130_fd_sc_hd__a21o_1
X_18499_ _02184_ _02196_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__xor2_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20530_ _03421_ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20461_ _03362_ _03363_ _03364_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__or3_1
XFILLER_193_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21013_ clknet_leaf_12_i_clk _00782_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11530_ _04244_ _04281_ _04289_ _04309_ _04140_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__a311o_1
XFILLER_11_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20728_ clknet_leaf_83_i_clk _00497_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11461_ _04142_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__clkbuf_8
XFILLER_17_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20659_ clknet_leaf_63_i_clk _00443_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-12\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13200_ _05930_ _05933_ _05936_ _05871_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__a31o_1
X_10412_ _03537_ vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11392_ rbzero.row_render.size\[6\] gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04172_
+ sky130_fd_sc_hd__or2_1
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14180_ _06914_ _06916_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__nand2_1
XFILLER_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13131_ _05867_ _05697_ _05688_ _05783_ _05826_ _05801_ vssd1 vssd1 vccd1 vccd1 _05868_
+ sky130_fd_sc_hd__mux4_1
X_10343_ _03501_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13062_ _05794_ _05798_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__nand2_1
XFILLER_140_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12013_ rbzero.tex_b1\[43\] rbzero.tex_b1\[42\] _04392_ vssd1 vssd1 vccd1 vccd1 _04788_
+ sky130_fd_sc_hd__mux2_1
X_17870_ _01471_ _01489_ _01487_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a21o_1
XFILLER_61_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16821_ _09461_ _09462_ vssd1 vssd1 vccd1 vccd1 _09463_ sky130_fd_sc_hd__or2_1
XFILLER_4_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16752_ _09254_ _09255_ vssd1 vssd1 vccd1 vccd1 _09394_ sky130_fd_sc_hd__or2_1
X_19540_ _03002_ _03000_ _03011_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__or3_1
X_13964_ _06696_ _06690_ _06672_ _06698_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__o22ai_1
XFILLER_4_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15703_ _08345_ _08346_ vssd1 vssd1 vccd1 vccd1 _08348_ sky130_fd_sc_hd__nor2_1
XFILLER_46_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12915_ _04031_ _05372_ _05651_ _04001_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__03040_ clknet_0__03040_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03040_
+ sky130_fd_sc_hd__clkbuf_16
X_16683_ _09186_ _09187_ _09325_ vssd1 vssd1 vccd1 vccd1 _09326_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19471_ rbzero.wall_tracer.rayAddendY\[4\] rbzero.wall_tracer.rayAddendY\[3\] _02904_
+ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__o21ai_2
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13895_ _06620_ _06631_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__or2_1
XFILLER_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18422_ _02118_ _02119_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__nand2_1
X_15634_ _08252_ _08261_ vssd1 vssd1 vccd1 vccd1 _08279_ sky130_fd_sc_hd__nor2_1
XFILLER_62_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12846_ rbzero.wall_tracer.visualWallDist\[-7\] _05351_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__mux2_1
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _02049_ _02051_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__xor2_1
XFILLER_15_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15565_ _08208_ _08209_ _05194_ vssd1 vssd1 vccd1 vccd1 _08210_ sky130_fd_sc_hd__o21ai_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12777_ _05519_ _05521_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _09864_ _09866_ _09865_ vssd1 vssd1 vccd1 vccd1 _09875_ sky130_fd_sc_hd__a21boi_1
XFILLER_202_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14516_ _07067_ _07069_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__nor2_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18284_ _01982_ _01983_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ rbzero.debug_overlay.playerY\[-7\] _04455_ _04501_ _04504_ _04506_ vssd1
+ vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a2111o_1
X_15496_ _08097_ _08128_ vssd1 vssd1 vccd1 vccd1 _08141_ sky130_fd_sc_hd__or2_1
X_17235_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _09813_ sky130_fd_sc_hd__or2_1
X_14447_ _07168_ _07183_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11659_ _04424_ _04426_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__nor2_1
XFILLER_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17166_ rbzero.traced_texa\[-4\] _09768_ _09767_ rbzero.wall_tracer.visualWallDist\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__a22o_1
XFILLER_196_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14378_ _06724_ _06740_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__or2_1
XFILLER_155_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16117_ _08739_ _08760_ vssd1 vssd1 vccd1 vccd1 _08762_ sky130_fd_sc_hd__nor2_1
X_13329_ _05752_ _06053_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__nand2_1
X_17097_ _09735_ _09736_ vssd1 vssd1 vccd1 vccd1 _09737_ sky130_fd_sc_hd__nor2_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20252__271 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__inv_2
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16048_ _08654_ _08663_ vssd1 vssd1 vccd1 vccd1 _08693_ sky130_fd_sc_hd__xnor2_2
XFILLER_171_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19628__80 clknet_1_0__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__inv_2
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19807_ _03132_ vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17999_ _09526_ _09480_ _09484_ _09391_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__o22a_1
XFILLER_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03307_ clknet_0__03307_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03307_
+ sky130_fd_sc_hd__clkbuf_16
X_19738_ rbzero.pov.spi_buffer\[43\] rbzero.pov.spi_buffer\[44\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03097_ sky130_fd_sc_hd__mux2_1
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19669_ rbzero.pov.spi_buffer\[10\] rbzero.pov.spi_buffer\[11\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03061_ sky130_fd_sc_hd__mux2_1
XFILLER_198_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21631_ clknet_leaf_29_i_clk _01400_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21562_ net483 _01331_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20513_ _03407_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__and2b_1
X_21493_ net414 _01262_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20335__346 clknet_1_1__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__inv_2
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20444_ rbzero.texV\[-7\] _03175_ _03332_ _03350_ vssd1 vssd1 vccd1 vccd1 _01389_
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20381__388 clknet_1_1__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__inv_2
XFILLER_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10961_ _03481_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__clkbuf_4
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12700_ rbzero.wall_tracer.rayAddendX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__or2_1
X_20080__116 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__inv_2
XFILLER_189_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13680_ _06395_ _06415_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__or2_1
X_10892_ rbzero.tex_b1\[44\] rbzero.tex_b1\[45\] _03784_ vssd1 vssd1 vccd1 vccd1 _03792_
+ sky130_fd_sc_hd__mux2_1
XFILLER_203_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12631_ rbzero.map_rom.d6 _05377_ _05375_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__a21oi_1
XFILLER_93_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15350_ _07990_ rbzero.wall_tracer.stepDistX\[-3\] _07994_ vssd1 vssd1 vccd1 vccd1
+ _07995_ sky130_fd_sc_hd__o21bai_4
XFILLER_157_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12562_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__nor2_1
XFILLER_157_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14301_ _07034_ _07036_ _07037_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__and3_1
X_11513_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _04291_ vssd1 vssd1 vccd1 vccd1 _04293_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15281_ _05346_ _05468_ _07893_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__mux2_1
XFILLER_184_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12493_ rbzero.wall_tracer.trackDistY\[-7\] _05238_ _05239_ rbzero.wall_tracer.trackDistY\[-8\]
+ _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__o221a_1
XFILLER_200_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17020_ _09539_ _09548_ _09547_ vssd1 vssd1 vccd1 vccd1 _09660_ sky130_fd_sc_hd__a21o_2
XFILLER_184_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14232_ _06942_ _06943_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__or2_1
X_11444_ _04138_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__buf_4
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _06893_ _06898_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__nor2_1
X_11375_ rbzero.row_render.size\[7\] rbzero.row_render.size\[6\] rbzero.row_render.size\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__a21o_1
XFILLER_3_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13114_ _05820_ _05849_ _05850_ _05798_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__o211a_1
XFILLER_180_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10326_ _03492_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14094_ _06827_ _06829_ _06830_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__a21oi_1
X_18971_ _02615_ vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _09103_ _09552_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__or2_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _05781_ _05702_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__or2_1
XFILLER_191_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17853_ _10179_ _10181_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__or2_1
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16804_ _09309_ _09311_ vssd1 vssd1 vccd1 vccd1 _09446_ sky130_fd_sc_hd__and2_1
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17784_ _01485_ _01486_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__and2_1
XFILLER_66_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14996_ _07668_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19523_ _02979_ _02989_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__or2_1
X_16735_ _09375_ _09376_ vssd1 vssd1 vccd1 vccd1 _09377_ sky130_fd_sc_hd__nor2_1
X_13947_ _06673_ _06683_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16666_ _09305_ _09306_ _09308_ vssd1 vssd1 vccd1 vccd1 _09309_ sky130_fd_sc_hd__nand3_1
X_19454_ _02923_ _02925_ _02935_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__or3_1
X_13878_ _06598_ _06599_ _06614_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__a21oi_4
XFILLER_90_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18405_ _01966_ _02000_ _02103_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__a21oi_2
X_15617_ _08252_ _08261_ vssd1 vssd1 vccd1 vccd1 _08262_ sky130_fd_sc_hd__xor2_1
XFILLER_201_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12829_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__buf_2
X_16597_ _09098_ _09108_ _09106_ vssd1 vssd1 vccd1 vccd1 _09240_ sky130_fd_sc_hd__a21o_1
X_19385_ _02870_ _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18336_ _01987_ _01994_ _02034_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__a21o_1
X_15548_ _08179_ _08190_ _08192_ vssd1 vssd1 vccd1 vccd1 _08193_ sky130_fd_sc_hd__a21o_1
XFILLER_203_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18267_ _08895_ _08767_ _01524_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__or3_1
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15479_ _07951_ _08123_ _08062_ _05207_ vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__a211o_4
XFILLER_147_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17218_ _09792_ _09796_ _09797_ vssd1 vssd1 vccd1 vccd1 _09799_ sky130_fd_sc_hd__o21ai_1
X_18198_ _01697_ _01780_ _01898_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a21oi_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17149_ rbzero.row_render.texu\[0\] _09762_ _07728_ rbzero.wall_tracer.texu\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__a22o_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20160_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__buf_1
XFILLER_116_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20993_ clknet_leaf_14_i_clk _00762_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_53_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21614_ clknet_leaf_35_i_clk _01383_ vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_205_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21545_ net466 _01314_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21476_ net397 _01245_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20427_ _03333_ _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03043_ clknet_0__03043_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03043_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11160_ rbzero.wall_tracer.mapX\[8\] _03947_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_
+ sky130_fd_sc_hd__or3b_1
XFILLER_1_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11091_ rbzero.tex_b0\[14\] rbzero.tex_b0\[13\] _03887_ vssd1 vssd1 vccd1 vccd1 _03896_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19607__61 clknet_1_1__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__inv_2
XFILLER_103_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14850_ _07569_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19622__75 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__inv_2
X_13801_ _05824_ _06535_ _06536_ _06537_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__or4_1
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14781_ _07487_ _07456_ _07513_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__a21oi_4
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11993_ rbzero.tex_b1\[1\] rbzero.tex_b1\[0\] _04250_ vssd1 vssd1 vccd1 vccd1 _04768_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16520_ _09163_ vssd1 vssd1 vccd1 vccd1 _09164_ sky130_fd_sc_hd__buf_2
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13732_ _06057_ _06045_ _05945_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__or3_1
XFILLER_204_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10944_ _03819_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16451_ _08821_ _08059_ _09094_ vssd1 vssd1 vccd1 vccd1 _09095_ sky130_fd_sc_hd__or3_1
XFILLER_43_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13663_ _06357_ _06399_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10875_ rbzero.tex_b1\[52\] rbzero.tex_b1\[53\] _03773_ vssd1 vssd1 vccd1 vccd1 _03783_
+ sky130_fd_sc_hd__mux2_1
X_15402_ _08046_ vssd1 vssd1 vccd1 vccd1 _08047_ sky130_fd_sc_hd__buf_4
XFILLER_25_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ gpout0.vpos\[9\] _04315_ _02703_ _02706_ vssd1 vssd1 vccd1 vccd1 _02727_
+ sky130_fd_sc_hd__or4_4
X_12614_ _05315_ _05366_ _05314_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__or3_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16382_ rbzero.wall_tracer.visualWallDist\[6\] _08148_ vssd1 vssd1 vccd1 vccd1 _09027_
+ sky130_fd_sc_hd__nand2_8
X_13594_ _06302_ _06329_ _06330_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__o21ba_1
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _01462_ _09480_ _09484_ _09526_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__o22a_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ rbzero.wall_tracer.visualWallDist\[-9\] _07903_ vssd1 vssd1 vccd1 vccd1 _07978_
+ sky130_fd_sc_hd__or2_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12545_ _05297_ _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__and2_1
XFILLER_184_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20318__330 clknet_1_0__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__inv_2
XFILLER_177_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18052_ _10125_ _10136_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__nand2_1
XFILLER_8_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15264_ _07908_ rbzero.debug_overlay.playerY\[-6\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _07909_ sky130_fd_sc_hd__mux2_1
XFILLER_200_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12476_ _05214_ rbzero.wall_tracer.trackDistX\[10\] _05230_ vssd1 vssd1 vccd1 vccd1
+ _05231_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17003_ _07994_ _08705_ _08058_ _08150_ vssd1 vssd1 vccd1 vccd1 _09643_ sky130_fd_sc_hd__or4_1
XFILLER_126_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14215_ _06852_ _06950_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__and2b_1
X_11427_ _04143_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__buf_6
XANTENNA_5 _05893_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _07820_ _07730_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__and2_1
XFILLER_99_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14146_ _06842_ _06881_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__and2_1
XFILLER_152_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11358_ _04089_ _04114_ _04124_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__nor3b_2
XFILLER_141_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10309_ rbzero.tex_r1\[63\] net46 _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__mux2_1
XFILLER_113_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14077_ _06800_ _06813_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__xnor2_1
X_18954_ rbzero.pov.spi_buffer\[10\] rbzero.pov.ready_buffer\[10\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02607_ sky130_fd_sc_hd__mux2_1
XFILLER_141_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11289_ _04065_ _04068_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__nor2_1
X_17905_ _01575_ _01607_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__xor2_1
X_13028_ _05567_ _05575_ _05656_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__o21a_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18885_ rbzero.spi_registers.new_vinf rbzero.spi_registers.spi_buffer\[0\] _02555_
+ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__mux2_1
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17836_ _10277_ _10279_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__or2b_1
XFILLER_67_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20364__372 clknet_1_0__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__inv_2
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17767_ _01461_ _01470_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__xor2_1
XFILLER_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14979_ _07659_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__clkbuf_1
X_20063__100 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__inv_2
X_19506_ _02963_ _02966_ _02964_ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a21boi_1
X_16718_ _08162_ _09214_ _09359_ _09212_ vssd1 vssd1 vccd1 vccd1 _09360_ sky130_fd_sc_hd__o31a_1
X_17698_ _10258_ _10262_ vssd1 vssd1 vccd1 vccd1 _10263_ sky130_fd_sc_hd__xor2_2
XFILLER_23_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19437_ _02920_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__clkbuf_1
X_16649_ _09288_ vssd1 vssd1 vccd1 vccd1 _09292_ sky130_fd_sc_hd__buf_4
XFILLER_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03037_ _03037_ vssd1 vssd1 vccd1 vccd1 clknet_0__03037_ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19368_ _07676_ _02856_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__nor2_1
XFILLER_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18319_ _01909_ _01911_ _01910_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__o21bai_1
XFILLER_202_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19299_ _02805_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21330_ net251 _01099_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21261_ clknet_leaf_96_i_clk _01030_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-5\]
+ sky130_fd_sc_hd__dfxtp_4
X_21192_ clknet_leaf_77_i_clk _00961_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20976_ clknet_leaf_8_i_clk _00745_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10660_ _03670_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10591_ _03633_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12330_ net29 _05089_ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__o21a_1
X_20192__217 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__inv_2
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21528_ net449 _01297_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12261_ net21 net22 _05027_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__and4_1
XFILLER_108_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21459_ net380 _01228_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14000_ _06735_ _06736_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__nor2_1
X_11212_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__buf_2
XFILLER_108_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12192_ _04960_ _04961_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__nor2_1
XFILLER_190_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput53 net53 vssd1 vssd1 vccd1 vccd1 o_gpout[0] sky130_fd_sc_hd__clkbuf_1
X_11143_ rbzero.debug_overlay.playerX\[2\] _03929_ rbzero.map_rom.d6 _03930_ _03931_
+ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__a221o_1
XFILLER_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput64 net64 vssd1 vssd1 vccd1 vccd1 o_rgb[23] sky130_fd_sc_hd__buf_2
XFILLER_123_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11074_ _03717_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__clkbuf_4
X_15951_ _08591_ _08592_ vssd1 vssd1 vccd1 vccd1 _08596_ sky130_fd_sc_hd__nand2_1
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14902_ _07591_ _07608_ _07609_ _04039_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__o211a_1
X_18670_ _08445_ _09704_ _02256_ _02365_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__o31a_1
X_15882_ _08476_ _08473_ vssd1 vssd1 vccd1 vccd1 _08527_ sky130_fd_sc_hd__nand2_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ _09912_ _10047_ _10045_ vssd1 vssd1 vccd1 vccd1 _10186_ sky130_fd_sc_hd__a21o_1
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ _07459_ _07439_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__nor2_1
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ _10116_ _10117_ vssd1 vssd1 vccd1 vccd1 _10118_ sky130_fd_sc_hd__xnor2_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _07420_ _07347_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__nand2_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11976_ rbzero.tex_b1\[30\] _04272_ _04265_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a21o_1
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16503_ _08976_ _08990_ _09146_ vssd1 vssd1 vccd1 vccd1 _09147_ sky130_fd_sc_hd__a21oi_2
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13715_ _06441_ _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__or2_1
X_17483_ _09947_ _09949_ vssd1 vssd1 vccd1 vccd1 _10049_ sky130_fd_sc_hd__nor2_1
XFILLER_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10927_ _03810_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14695_ _07418_ _07422_ _07424_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__or4b_1
XFILLER_147_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19222_ rbzero.color_floor\[5\] _02751_ _02760_ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__a21o_1
X_13646_ _06382_ _05923_ _06116_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__and3_1
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16434_ _09077_ _09078_ vssd1 vssd1 vccd1 vccd1 _09079_ sky130_fd_sc_hd__nand2_1
X_10858_ _03774_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16365_ _07995_ _08109_ _08084_ _07931_ vssd1 vssd1 vccd1 vccd1 _09010_ sky130_fd_sc_hd__o22a_1
X_19153_ rbzero.spi_registers.new_other\[9\] _02712_ vssd1 vssd1 vccd1 vccd1 _02717_
+ sky130_fd_sc_hd__or2_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13577_ _06312_ _06313_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__xnor2_1
X_10789_ rbzero.tex_g0\[30\] rbzero.tex_g0\[29\] _03729_ vssd1 vssd1 vccd1 vccd1 _03738_
+ sky130_fd_sc_hd__mux2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18104_ _01700_ _01731_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__or2_1
XFILLER_200_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15316_ rbzero.wall_tracer.state\[3\] _07960_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__nand2_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12528_ _05203_ _05211_ _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__o21ai_4
X_19084_ _02674_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__clkbuf_1
X_16296_ _08719_ _08763_ vssd1 vssd1 vccd1 vccd1 _08941_ sky130_fd_sc_hd__nor2_1
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18035_ _08493_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__buf_2
X_15247_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__clkbuf_4
X_12459_ rbzero.wall_tracer.trackDistY\[10\] vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__inv_2
XFILLER_114_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15178_ _07816_ _07824_ _07828_ _07831_ vssd1 vssd1 vccd1 vccd1 _07832_ sky130_fd_sc_hd__a31o_1
XFILLER_158_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14129_ _06769_ _06662_ _06667_ _06776_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__o22a_1
XFILLER_141_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19986_ _02721_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18937_ rbzero.pov.spi_buffer\[2\] rbzero.pov.ready_buffer\[2\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02598_ sky130_fd_sc_hd__mux2_1
XFILLER_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18868_ _02540_ _02541_ _02228_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__o21ai_1
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17819_ _01516_ _01522_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__xor2_1
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18799_ _02479_ _02476_ _02480_ _02481_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__a211o_1
XFILLER_36_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20830_ clknet_leaf_51_i_clk _00599_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19601__56 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__inv_2
XFILLER_63_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20761_ clknet_leaf_46_i_clk _00530_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20692_ clknet_leaf_57_i_clk _00476_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21313_ net234 _01082_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21244_ clknet_leaf_91_i_clk _01013_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21175_ clknet_leaf_5_i_clk _00944_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ rbzero.tex_g1\[59\] rbzero.tex_g1\[58\] _04337_ vssd1 vssd1 vccd1 vccd1 _04607_
+ sky130_fd_sc_hd__mux2_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _04119_ _04526_ _04530_ _04538_ _04121_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__o311a_1
X_20959_ clknet_leaf_1_i_clk _00728_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13500_ _06160_ _06202_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__nand2_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _03697_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14480_ _07200_ _07215_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__nor2_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ rbzero.debug_overlay.vplaneY\[-3\] vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__buf_4
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20200__224 clknet_1_0__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__inv_2
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _06156_ _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__nor2_1
X_10643_ _03661_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16150_ _08780_ _08781_ vssd1 vssd1 vccd1 vccd1 _08795_ sky130_fd_sc_hd__nand2_1
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13362_ _06025_ _06027_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10574_ rbzero.tex_r0\[4\] rbzero.tex_r0\[3\] _03624_ vssd1 vssd1 vccd1 vccd1 _03625_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15101_ _07741_ _07744_ vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__or2_1
X_12313_ net30 net31 vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__nor2_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16081_ _08723_ _08724_ vssd1 vssd1 vccd1 vccd1 _08726_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13293_ _06024_ _06028_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__xor2_1
XFILLER_138_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15032_ rbzero.debug_overlay.vplaneX\[-9\] _03914_ _07679_ _07694_ _07696_ vssd1
+ vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__a221o_1
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12244_ net48 net39 net38 net40 net15 _04961_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__mux4_1
XFILLER_6_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19840_ _03139_ _03154_ _03156_ _03157_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__o211a_1
X_12175_ _04892_ _04909_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__o21a_1
XFILLER_123_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11126_ rbzero.wall_tracer.visualWallDist\[0\] rbzero.wall_tracer.visualWallDist\[-1\]
+ rbzero.wall_tracer.visualWallDist\[-2\] rbzero.wall_tracer.visualWallDist\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__or4_1
XFILLER_95_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19771_ _03046_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__buf_4
XFILLER_68_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16983_ _08331_ _09621_ _09488_ _09622_ vssd1 vssd1 vccd1 vccd1 _09623_ sky130_fd_sc_hd__a31oi_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20407__8 clknet_1_1__leaf__03037_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__inv_2
X_18722_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.stepDistY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__or2_1
XFILLER_95_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15934_ _08572_ vssd1 vssd1 vccd1 vccd1 _08579_ sky130_fd_sc_hd__buf_2
X_11057_ _03878_ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18653_ _02331_ _02348_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__xnor2_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ _08467_ _08464_ vssd1 vssd1 vccd1 vccd1 _08510_ sky130_fd_sc_hd__and2b_1
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _09906_ _10168_ _10169_ vssd1 vssd1 vccd1 vccd1 _10170_ sky130_fd_sc_hd__o21a_1
X_14816_ _07486_ _07399_ _07543_ _07527_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__a22o_1
X_18584_ _02271_ _02280_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__xnor2_1
Xtop_ew_algofoogle_110 vssd1 vssd1 vccd1 vccd1 ones[4] top_ew_algofoogle_110/LO sky130_fd_sc_hd__conb_1
XFILLER_188_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _08391_ _08397_ vssd1 vssd1 vccd1 vccd1 _08441_ sky130_fd_sc_hd__xnor2_1
Xtop_ew_algofoogle_121 vssd1 vssd1 vccd1 vccd1 ones[15] top_ew_algofoogle_121/LO sky130_fd_sc_hd__conb_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17535_ _09670_ _10099_ _10100_ vssd1 vssd1 vccd1 vccd1 _10101_ sky130_fd_sc_hd__a21o_1
XFILLER_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11959_ _04206_ _04700_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__and3b_1
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14747_ _07473_ _07478_ _07481_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__o21bai_1
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14678_ _07378_ _07413_ _07414_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__nor3_1
X_17466_ _10032_ vssd1 vssd1 vccd1 vccd1 _10033_ sky130_fd_sc_hd__inv_2
XFILLER_189_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19205_ _09753_ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__and2_1
X_13629_ _06355_ _06359_ _06365_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__o21ba_1
X_16417_ _08549_ _08957_ _09060_ vssd1 vssd1 vccd1 vccd1 _09062_ sky130_fd_sc_hd__nand3_4
XFILLER_32_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17397_ _09126_ _08570_ vssd1 vssd1 vccd1 vccd1 _09964_ sky130_fd_sc_hd__nor2_1
XFILLER_34_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20175__201 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__inv_2
XFILLER_186_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19136_ _04891_ _04887_ gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__nand3_2
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16348_ _08206_ _08248_ _08992_ vssd1 vssd1 vccd1 vccd1 _08993_ sky130_fd_sc_hd__a21o_1
X_16279_ _08876_ _08923_ vssd1 vssd1 vccd1 vccd1 _08924_ sky130_fd_sc_hd__nand2_1
X_19067_ rbzero.pov.spi_buffer\[64\] rbzero.pov.ready_buffer\[64\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02666_ sky130_fd_sc_hd__mux2_1
XFILLER_173_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18018_ _01718_ _01719_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__nand2_1
XFILLER_161_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19969_ rbzero.pov.ready_buffer\[42\] _03240_ _03243_ rbzero.debug_overlay.facingX\[0\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__o221a_1
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20813_ clknet_leaf_55_i_clk _00582_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20744_ clknet_leaf_43_i_clk _00513_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20675_ clknet_leaf_48_i_clk _00459_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_104_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03291_ clknet_0__03291_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03291_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21227_ clknet_leaf_21_i_clk _00996_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_137_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21158_ clknet_leaf_68_i_clk _00927_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13980_ _06245_ _06678_ _06715_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__o21bai_1
X_21089_ net179 _00858_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12931_ _05628_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__nand2_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15650_ _08289_ _08294_ vssd1 vssd1 vccd1 vccd1 _08295_ sky130_fd_sc_hd__xnor2_2
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _05594_ _05596_ _05598_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__nor3_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _04205_ _04556_ _04590_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__and3b_1
X_14601_ _07327_ _07326_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__and2b_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ rbzero.wall_tracer.visualWallDist\[-11\] _04012_ vssd1 vssd1 vccd1 vccd1
+ _08226_ sky130_fd_sc_hd__nand2_4
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ rbzero.wall_tracer.mapY\[5\] _05397_ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_
+ sky130_fd_sc_hd__o21a_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14532_ _07254_ _07257_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__nand2_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _05394_ vssd1 vssd1 vccd1 vccd1 _09889_ sky130_fd_sc_hd__clkbuf_4
XFILLER_183_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11744_ _04522_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_8
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _07160_ _07199_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__nor2_1
X_17251_ _09824_ _09825_ _09827_ vssd1 vssd1 vccd1 vccd1 _09828_ sky130_fd_sc_hd__o21ai_1
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11675_ _04433_ _04447_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__and2_2
XFILLER_186_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16202_ _08840_ _08846_ vssd1 vssd1 vccd1 vccd1 _08847_ sky130_fd_sc_hd__nand2_1
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ _06021_ _06050_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__and2b_1
X_10626_ _03652_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__clkbuf_1
X_17182_ rbzero.traced_texa\[9\] _09770_ _09771_ rbzero.wall_tracer.visualWallDist\[9\]
+ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__a22o_1
X_14394_ _07111_ _07128_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__nand2_1
X_16133_ _08660_ _08777_ vssd1 vssd1 vccd1 vccd1 _08778_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ _06063_ _06081_ _06073_ _06070_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__a2bb2o_1
X_10557_ rbzero.tex_r0\[12\] rbzero.tex_r0\[11\] _03613_ vssd1 vssd1 vccd1 vccd1 _03616_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16064_ _08701_ _08708_ vssd1 vssd1 vccd1 vccd1 _08709_ sky130_fd_sc_hd__xor2_2
X_13276_ _05978_ _05981_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__nor2_1
X_10488_ _03579_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15015_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.wall_tracer.rayAddendX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__nor2_1
XFILLER_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12227_ net49 _04962_ _04980_ net52 vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a22o_1
XFILLER_190_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20170__197 clknet_1_1__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__inv_2
X_19823_ _03139_ _03142_ _03144_ _02765_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__o211a_1
XFILLER_97_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12158_ _04323_ _04903_ _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a21o_1
XFILLER_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11109_ _03905_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__clkbuf_1
X_19754_ _03105_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12089_ _04858_ _04860_ net5 vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__mux2_1
X_16966_ _09345_ _09590_ vssd1 vssd1 vccd1 vccd1 _09606_ sky130_fd_sc_hd__and2_1
X_18705_ rbzero.wall_tracer.trackDistY\[-12\] _02397_ _02399_ vssd1 vssd1 vccd1 vccd1
+ _02400_ sky130_fd_sc_hd__mux2_1
X_15917_ _08482_ _08559_ _08560_ _08561_ vssd1 vssd1 vccd1 vccd1 _08562_ sky130_fd_sc_hd__a2bb2o_1
X_19685_ rbzero.pov.spi_buffer\[18\] rbzero.pov.spi_buffer\[19\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03069_ sky130_fd_sc_hd__mux2_1
X_16897_ _09518_ _09537_ vssd1 vssd1 vccd1 vccd1 _09538_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18636_ _02273_ _02274_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__and2_1
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _08129_ vssd1 vssd1 vccd1 vccd1 _08493_ sky130_fd_sc_hd__buf_4
XFILLER_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18567_ _01498_ _09215_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__nor2_1
XFILLER_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15779_ _05208_ _08423_ vssd1 vssd1 vccd1 vccd1 _08424_ sky130_fd_sc_hd__or2_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17518_ _10069_ _10083_ vssd1 vssd1 vccd1 vccd1 _10084_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18498_ _02193_ _02195_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__xor2_1
XFILLER_33_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17449_ _09722_ _09724_ vssd1 vssd1 vccd1 vccd1 _10016_ sky130_fd_sc_hd__nor2_1
XFILLER_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20460_ _03357_ _03359_ _03358_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__a21boi_1
XFILLER_192_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19119_ rbzero.spi_registers.spi_cmd\[2\] rbzero.spi_registers.spi_cmd\[3\] _02690_
+ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__mux2_1
XFILLER_145_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21012_ clknet_leaf_12_i_clk _00781_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20147__177 clknet_1_1__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__inv_2
XFILLER_43_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20727_ clknet_leaf_80_i_clk _00496_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ _04237_ _04238_ _04239_ _04226_ _04210_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__o221a_1
XFILLER_184_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20658_ clknet_leaf_51_i_clk _00442_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_139_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10411_ rbzero.tex_r1\[14\] rbzero.tex_r1\[15\] _03527_ vssd1 vssd1 vccd1 vccd1 _03537_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11391_ rbzero.row_render.size\[6\] gpout0.hpos\[6\] _04004_ _04160_ _04170_ vssd1
+ vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__a221o_1
X_20589_ _03456_ _03457_ rbzero.wall_tracer.rayAddendX\[-6\] _09762_ vssd1 vssd1 vccd1
+ vccd1 _01427_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_178_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13130_ _05710_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__inv_2
X_10342_ rbzero.tex_r1\[47\] rbzero.tex_r1\[48\] _03494_ vssd1 vssd1 vccd1 vccd1 _03501_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20312__325 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__inv_2
XFILLER_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _05754_ _05797_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__nand2_2
XFILLER_151_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12012_ _04242_ _04778_ _04786_ _04207_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__o211a_1
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16820_ _09458_ _09460_ vssd1 vssd1 vccd1 vccd1 _09462_ sky130_fd_sc_hd__and2_1
XFILLER_120_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16751_ _09390_ _09392_ vssd1 vssd1 vccd1 vccd1 _09393_ sky130_fd_sc_hd__and2_1
XFILLER_120_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13963_ _06697_ _06699_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__nand2_2
XFILLER_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15702_ _08345_ _08346_ vssd1 vssd1 vccd1 vccd1 _08347_ sky130_fd_sc_hd__xor2_1
XFILLER_47_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19470_ _02925_ _02935_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__nand2_1
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12914_ rbzero.wall_tracer.visualWallDist\[6\] _04031_ vssd1 vssd1 vccd1 vccd1 _05651_
+ sky130_fd_sc_hd__nor2_1
X_16682_ _09183_ _09185_ vssd1 vssd1 vccd1 vccd1 _09325_ sky130_fd_sc_hd__or2_1
XFILLER_46_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13894_ _06629_ _06630_ vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__nand2_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18421_ _02118_ _02119_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__or2_1
XFILLER_59_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15633_ _08268_ _08277_ vssd1 vssd1 vccd1 vccd1 _08278_ sky130_fd_sc_hd__xnor2_1
X_12845_ _05561_ _05469_ _05580_ _05581_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__o22a_2
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18352_ _10248_ _09977_ _01990_ _02050_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__o31a_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _05513_ _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__nand2_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _07560_ _07562_ _08171_ _07564_ vssd1 vssd1 vccd1 vccd1 _08209_ sky130_fd_sc_hd__o31a_1
XFILLER_199_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _09872_ _09873_ vssd1 vssd1 vccd1 vccd1 _09874_ sky130_fd_sc_hd__or2b_1
X_14515_ _07235_ _07251_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__xnor2_1
X_11727_ rbzero.debug_overlay.playerY\[3\] _04452_ _04464_ rbzero.debug_overlay.playerY\[-4\]
+ _04505_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__a221o_1
X_18283_ _09141_ _10238_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__nor2_1
X_15495_ _08109_ _08104_ _08042_ _08084_ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__o22a_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17234_ _04016_ vssd1 vssd1 vccd1 vccd1 _09812_ sky130_fd_sc_hd__buf_4
XFILLER_31_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14446_ _07170_ _07182_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__xor2_1
X_11658_ _04422_ _04436_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__nor2_1
X_10609_ rbzero.tex_g1\[50\] rbzero.tex_g1\[51\] _03635_ vssd1 vssd1 vccd1 vccd1 _03643_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14377_ _07112_ _07113_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__nor2_1
X_17165_ rbzero.traced_texa\[-5\] _09768_ _09767_ rbzero.wall_tracer.visualWallDist\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__a22o_1
X_11589_ rbzero.tex_r1\[31\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__and3_1
XFILLER_122_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13328_ _05852_ _05853_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__nand2_4
X_16116_ _08739_ _08760_ vssd1 vssd1 vccd1 vccd1 _08761_ sky130_fd_sc_hd__xor2_2
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17096_ _09605_ _09606_ _09734_ vssd1 vssd1 vccd1 vccd1 _09736_ sky130_fd_sc_hd__o21a_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13259_ _05988_ _05989_ _05992_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__a22o_1
X_16047_ _08682_ _08689_ _08691_ vssd1 vssd1 vccd1 vccd1 _08692_ sky130_fd_sc_hd__a21oi_4
XFILLER_170_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20287__302 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__inv_2
XFILLER_142_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19806_ rbzero.pov.ss_buffer\[1\] rbzero.pov.ss_buffer\[0\] _05189_ vssd1 vssd1 vccd1
+ vccd1 _03132_ sky130_fd_sc_hd__mux2_1
X_17998_ _01613_ _01631_ _01699_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03306_ clknet_0__03306_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03306_
+ sky130_fd_sc_hd__clkbuf_16
X_19737_ _03096_ vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__clkbuf_1
X_16949_ _09587_ _09589_ vssd1 vssd1 vccd1 vccd1 _09590_ sky130_fd_sc_hd__xor2_1
XFILLER_84_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20402__27 clknet_1_1__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__inv_2
XFILLER_38_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19668_ _03060_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18619_ _02313_ _02315_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__or2_1
XFILLER_80_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21630_ clknet_leaf_31_i_clk _01399_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21561_ net482 _01330_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20512_ rbzero.traced_texa\[4\] rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _03408_
+ sky130_fd_sc_hd__nand2_1
X_21492_ net413 _01261_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20443_ _03348_ _03349_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_51_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_10_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_66_i_clk clknet_opt_13_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10960_ _03827_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10891_ _03791_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12630_ _05381_ _05382_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__nor2_1
XFILLER_58_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12561_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__and2_1
XFILLER_106_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11512_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _04291_ vssd1 vssd1 vccd1 vccd1 _04292_
+ sky130_fd_sc_hd__mux2_1
X_14300_ _06911_ _06914_ _06884_ _06885_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__a211oi_2
XFILLER_12_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15280_ _04013_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__clkbuf_8
XFILLER_200_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12492_ _05239_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.trackDistY\[-9\]
+ _05240_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__a221o_1
XFILLER_156_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ _06888_ _06966_ _06963_ _06940_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__o211ai_1
X_11443_ rbzero.tex_r0\[57\] _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__and3_1
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_184_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14162_ _06893_ _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__nand2_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11374_ gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13113_ _05797_ _05809_ _05839_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a21o_1
X_10325_ rbzero.tex_r1\[55\] rbzero.tex_r1\[56\] _03483_ vssd1 vssd1 vccd1 vccd1 _03492_
+ sky130_fd_sc_hd__mux2_1
X_14093_ _06804_ _06828_ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__and2b_1
X_18970_ rbzero.pov.spi_buffer\[18\] rbzero.pov.ready_buffer\[18\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02615_ sky130_fd_sc_hd__mux2_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _01503_ _01623_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13044_ _05695_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__clkinv_2
XFILLER_26_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17852_ _01554_ _01555_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__nand2_1
XFILLER_113_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16803_ _09405_ _09444_ vssd1 vssd1 vccd1 vccd1 _09445_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17783_ _01485_ _01486_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__nor2_1
XFILLER_207_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14995_ rbzero.wall_tracer.stepDistX\[4\] _07566_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07668_ sky130_fd_sc_hd__mux2_1
X_19522_ rbzero.wall_tracer.rayAddendY\[8\] _00013_ _02992_ _02999_ vssd1 vssd1 vccd1
+ vccd1 _00818_ sky130_fd_sc_hd__o22a_1
X_16734_ _09372_ _09374_ vssd1 vssd1 vccd1 vccd1 _09376_ sky130_fd_sc_hd__and2_1
X_13946_ _06674_ _06679_ _06682_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__a21oi_1
XFILLER_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20282__298 clknet_1_0__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__inv_2
XFILLER_62_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19453_ _02904_ rbzero.wall_tracer.rayAddendY\[4\] vssd1 vssd1 vccd1 vccd1 _02935_
+ sky130_fd_sc_hd__xor2_1
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16665_ _09125_ _09148_ _09307_ vssd1 vssd1 vccd1 vccd1 _09308_ sky130_fd_sc_hd__a21o_1
X_13877_ _06563_ _06600_ _06613_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__o21ai_2
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18404_ _01998_ _01999_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__nor2_1
X_15616_ _08256_ _08258_ _08260_ vssd1 vssd1 vccd1 vccd1 _08261_ sky130_fd_sc_hd__a21boi_1
X_19384_ _02860_ _02863_ _02861_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a21bo_1
X_12828_ _04030_ _05327_ _05371_ _05564_ _04001_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__a311o_1
X_16596_ _09209_ _09238_ vssd1 vssd1 vccd1 vccd1 _09239_ sky130_fd_sc_hd__xnor2_1
XFILLER_201_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18335_ _01992_ _01993_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__nor2_1
XFILLER_43_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15547_ _08170_ _08189_ _08191_ vssd1 vssd1 vccd1 vccd1 _08192_ sky130_fd_sc_hd__o21ba_1
XFILLER_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12759_ _05504_ _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__nor2_1
XFILLER_203_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18266_ _01929_ _01965_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__xnor2_2
XFILLER_129_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15478_ rbzero.wall_tracer.stepDistY\[-11\] vssd1 vssd1 vccd1 vccd1 _08123_ sky130_fd_sc_hd__inv_2
XFILLER_129_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17217_ _09792_ _09796_ _09797_ vssd1 vssd1 vccd1 vccd1 _09798_ sky130_fd_sc_hd__or3_1
X_14429_ _06696_ _06663_ _06708_ _06698_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__o22a_1
X_18197_ _01777_ _01779_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__nor2_1
XFILLER_157_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17148_ rbzero.row_render.size\[10\] _09762_ _07562_ _07756_ vssd1 vssd1 vccd1 vccd1
+ _00538_ sky130_fd_sc_hd__a22o_1
XFILLER_115_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17079_ _09571_ _09573_ vssd1 vssd1 vccd1 vccd1 _09719_ sky130_fd_sc_hd__and2b_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20992_ clknet_leaf_14_i_clk _00761_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20341__351 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__inv_2
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21613_ clknet_leaf_35_i_clk _01382_ vssd1 vssd1 vccd1 vccd1 gpout5.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21544_ net465 _01313_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20259__278 clknet_1_0__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__inv_2
XFILLER_166_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21475_ net396 _01244_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20426_ _03334_ _03335_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__and2b_1
XFILLER_101_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03042_ clknet_0__03042_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03042_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_146_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11090_ _03895_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ _06529_ _06533_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__nor2_1
XFILLER_21_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11992_ rbzero.tex_b1\[2\] _04272_ _04265_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__a21o_1
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14780_ _07459_ _07505_ _07510_ _07512_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__a31o_1
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13731_ _06448_ _06450_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__xor2_1
X_10943_ rbzero.tex_b1\[20\] rbzero.tex_b1\[21\] _03817_ vssd1 vssd1 vccd1 vccd1 _03819_
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16450_ _09092_ _09093_ vssd1 vssd1 vccd1 vccd1 _09094_ sky130_fd_sc_hd__nand2_1
X_10874_ _03782_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13662_ _06313_ _06356_ _06358_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__o21bai_1
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _08045_ vssd1 vssd1 vccd1 vccd1 _08046_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12613_ _05315_ _05366_ _05314_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__o21ai_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16381_ _08369_ _08349_ vssd1 vssd1 vccd1 vccd1 _09026_ sky130_fd_sc_hd__or2b_1
X_13593_ _06303_ _06328_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nor2_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _01735_ _01752_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a21oi_1
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12544_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__or2_1
X_15332_ _05208_ rbzero.wall_tracer.stepDistX\[-2\] _07976_ vssd1 vssd1 vccd1 vccd1
+ _07977_ sky130_fd_sc_hd__a21boi_4
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18051_ _01735_ _01752_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__xor2_1
XFILLER_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15263_ _07906_ _07907_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__and2_1
X_12475_ _05212_ rbzero.wall_tracer.trackDistY\[11\] vssd1 vssd1 vccd1 vccd1 _05230_
+ sky130_fd_sc_hd__nor2_1
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03309_ clknet_0__03309_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03309_
+ sky130_fd_sc_hd__clkbuf_16
X_17002_ _07994_ _08058_ _08151_ _08705_ vssd1 vssd1 vccd1 vccd1 _09642_ sky130_fd_sc_hd__o22a_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11426_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__clkbuf_4
X_14214_ _06950_ _06852_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__and2b_1
X_15194_ _07820_ _07730_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__nor2_1
XANTENNA_6 _07514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ _06842_ _06881_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__nor2_2
X_11357_ _04135_ _04136_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__and2_1
XFILLER_99_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ _03482_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__clkbuf_4
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14076_ _06802_ _06811_ _06812_ vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__a21oi_1
X_18953_ _02606_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11288_ rbzero.texV\[5\] _04066_ _04067_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__a21boi_1
X_17904_ _01591_ _01606_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__xnor2_1
X_13027_ _05574_ _05662_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__xor2_1
XFILLER_117_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18884_ rbzero.spi_registers.spi_done _03480_ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_
+ sky130_fd_sc_hd__and3_1
XFILLER_67_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17835_ _01492_ _01538_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17766_ _01468_ _01469_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__nor2_1
XFILLER_82_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14978_ rbzero.wall_tracer.stepDistX\[-4\] _07541_ _07650_ vssd1 vssd1 vccd1 vccd1
+ _07659_ sky130_fd_sc_hd__mux2_1
XFILLER_75_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19505_ _02982_ _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__nand2_1
X_16717_ _09217_ vssd1 vssd1 vccd1 vccd1 _09359_ sky130_fd_sc_hd__clkbuf_4
X_13929_ _05982_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__clkbuf_4
XFILLER_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17697_ _10260_ _10261_ vssd1 vssd1 vccd1 vccd1 _10262_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19436_ rbzero.wall_tracer.rayAddendY\[2\] _02919_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _02920_ sky130_fd_sc_hd__mux2_1
X_16648_ _08239_ _09288_ _09289_ _09290_ vssd1 vssd1 vccd1 vccd1 _09291_ sky130_fd_sc_hd__or4bb_1
XFILLER_204_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19367_ _02853_ _02855_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__xnor2_1
X_16579_ _09220_ _09221_ vssd1 vssd1 vccd1 vccd1 _09222_ sky130_fd_sc_hd__and2_1
XFILLER_124_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18318_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.stepDistX\[7\] vssd1
+ vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__nand2_1
XFILLER_198_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19298_ rbzero.spi_registers.new_other\[3\] rbzero.spi_registers.spi_buffer\[3\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__mux2_1
XFILLER_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18249_ _01938_ _01948_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__nand2_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21260_ clknet_leaf_88_i_clk _01029_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21191_ clknet_leaf_77_i_clk _00960_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20975_ clknet_leaf_15_i_clk _00744_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10590_ rbzero.tex_g1\[59\] rbzero.tex_g1\[60\] _03549_ vssd1 vssd1 vccd1 vccd1 _03633_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21527_ net448 _01296_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _05021_ net66 _05028_ net24 vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__a211o_1
XFILLER_107_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21458_ net379 _01227_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11211_ _03914_ _03999_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__nor2_1
X_20409_ gpout5.clk_div\[1\] gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__nand2_1
X_12191_ net14 vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__clkbuf_4
XFILLER_147_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21389_ net310 _01158_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11142_ rbzero.debug_overlay.playerY\[5\] rbzero.wall_tracer.mapY\[5\] vssd1 vssd1
+ vccd1 vccd1 _03931_ sky130_fd_sc_hd__xor2_1
Xoutput54 net510 vssd1 vssd1 vccd1 vccd1 o_gpout[1] sky130_fd_sc_hd__clkbuf_1
Xoutput65 net65 vssd1 vssd1 vccd1 vccd1 o_rgb[6] sky130_fd_sc_hd__buf_2
XFILLER_163_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11073_ _03886_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__clkbuf_1
X_15950_ _07974_ _08594_ vssd1 vssd1 vccd1 vccd1 _08595_ sky130_fd_sc_hd__or2_1
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14901_ rbzero.wall_tracer.visualWallDist\[-7\] _07595_ vssd1 vssd1 vccd1 vccd1 _07609_
+ sky130_fd_sc_hd__or2_1
XFILLER_114_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15881_ _08517_ _08525_ vssd1 vssd1 vccd1 vccd1 _08526_ sky130_fd_sc_hd__xor2_2
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17620_ _10169_ _10166_ _10165_ vssd1 vssd1 vccd1 vccd1 _10185_ sky130_fd_sc_hd__a21oi_1
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14832_ _00004_ _07555_ _07556_ vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__a21oi_1
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ _09114_ _09552_ vssd1 vssd1 vccd1 vccd1 _10117_ sky130_fd_sc_hd__nor2_1
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14763_ _07419_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__clkinv_2
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11975_ rbzero.tex_b1\[31\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__and3_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _08989_ _08987_ vssd1 vssd1 vccd1 vccd1 _09146_ sky130_fd_sc_hd__and2b_1
XFILLER_44_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13714_ _06442_ _06447_ _06448_ _06450_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17482_ _09912_ _10047_ vssd1 vssd1 vccd1 vccd1 _10048_ sky130_fd_sc_hd__xor2_1
X_10926_ rbzero.tex_b1\[28\] rbzero.tex_b1\[29\] _03806_ vssd1 vssd1 vccd1 vccd1 _03810_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14694_ _05742_ _07426_ _07430_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__a21o_1
XFILLER_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19221_ rbzero.spi_registers.new_floor\[5\] rbzero.spi_registers.got_new_floor _02711_
+ _03911_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__a31o_1
XFILLER_73_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16433_ _09074_ _09075_ vssd1 vssd1 vccd1 vccd1 _09078_ sky130_fd_sc_hd__or2_1
X_10857_ rbzero.tex_b1\[61\] rbzero.tex_b1\[62\] _03773_ vssd1 vssd1 vccd1 vccd1 _03774_
+ sky130_fd_sc_hd__mux2_1
X_13645_ _06065_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__inv_2
XFILLER_204_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19152_ rbzero.otherx\[2\] _02710_ _02716_ _02714_ vssd1 vssd1 vccd1 vccd1 _00731_
+ sky130_fd_sc_hd__o211a_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _07995_ _08570_ vssd1 vssd1 vccd1 vccd1 _09009_ sky130_fd_sc_hd__nor2_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10788_ _03737_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__clkbuf_1
X_13576_ _05946_ _05939_ _06007_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__or3_2
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _01563_ _01565_ _01696_ _01694_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__a31o_1
XFILLER_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15315_ _05360_ _05472_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__mux2_1
XFILLER_200_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19083_ rbzero.pov.spi_buffer\[72\] rbzero.pov.ready_buffer\[72\] _02594_ vssd1 vssd1
+ vccd1 vccd1 _02674_ sky130_fd_sc_hd__mux2_1
X_12527_ _04017_ _05279_ _05281_ _03970_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__o211a_1
X_16295_ _08851_ _08936_ _08937_ _08939_ vssd1 vssd1 vccd1 vccd1 _08940_ sky130_fd_sc_hd__o211a_1
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18034_ _01634_ _01642_ _01641_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a21bo_1
X_15246_ _07892_ vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__clkbuf_1
X_12458_ _05212_ rbzero.wall_tracer.trackDistY\[11\] vssd1 vssd1 vccd1 vccd1 _05213_
+ sky130_fd_sc_hd__and2_1
X_11409_ _04150_ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__nand2_1
X_12389_ net38 _05142_ _05139_ net48 _05155_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__a221o_1
XFILLER_125_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15177_ _07830_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__buf_6
XFILLER_207_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14128_ _06805_ _06707_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__or2_1
XFILLER_207_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19985_ rbzero.pov.ready_buffer\[12\] _03252_ _03253_ rbzero.debug_overlay.vplaneX\[-8\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__o221a_1
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14059_ _06786_ _06794_ _06795_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__a21bo_1
X_18936_ _02597_ vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_67_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18867_ _02537_ _02538_ _02539_ _04016_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__a31o_1
XFILLER_95_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19598__53 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__inv_2
X_17818_ _01517_ _01521_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__xor2_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18798_ _05257_ _08200_ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__nor2_1
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17749_ _01451_ _01452_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__nor2_1
XFILLER_36_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20760_ clknet_leaf_45_i_clk _00529_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_165_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19419_ _07756_ _02896_ _02897_ _02903_ vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__a31o_1
XFILLER_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20691_ clknet_leaf_58_i_clk _00475_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21312_ net233 _01081_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21243_ clknet_leaf_88_i_clk _01012_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_105_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21174_ clknet_leaf_6_i_clk _00943_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _04208_ _04533_ _04537_ _04142_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__a211o_1
XFILLER_198_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20958_ clknet_leaf_4_i_clk _00727_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ rbzero.tex_g1\[2\] rbzero.tex_g1\[3\] _03691_ vssd1 vssd1 vccd1 vccd1 _03697_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11691_ rbzero.debug_overlay.vplaneX\[10\] _04453_ _04457_ _04469_ vssd1 vssd1 vccd1
+ vccd1 _04470_ sky130_fd_sc_hd__a211o_1
XFILLER_42_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20889_ clknet_leaf_86_i_clk _00658_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10642_ rbzero.tex_g1\[35\] rbzero.tex_g1\[36\] _03658_ vssd1 vssd1 vccd1 vccd1 _03661_
+ sky130_fd_sc_hd__mux2_1
X_13430_ _06157_ _06166_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13361_ _06094_ _06095_ _06096_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__a21o_1
XFILLER_155_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10573_ _03557_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__clkbuf_4
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15100_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__or2_1
X_12312_ _05031_ _05041_ _05079_ _05080_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__o31a_2
XFILLER_182_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16080_ _08723_ _08724_ vssd1 vssd1 vccd1 vccd1 _08725_ sky130_fd_sc_hd__nand2_1
X_13292_ _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__inv_2
XFILLER_155_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12243_ net46 _04980_ _05012_ _05010_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__o2bb2a_1
X_15031_ rbzero.wall_tracer.rayAddendX\[-5\] _07695_ vssd1 vssd1 vccd1 vccd1 _07696_
+ sky130_fd_sc_hd__and2_1
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12174_ gpout0.vpos\[0\] net8 net10 net9 vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__o211a_1
XFILLER_190_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11125_ _03913_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__buf_4
X_19770_ _03113_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__clkbuf_1
X_16982_ _08329_ _09216_ _09351_ _08054_ vssd1 vssd1 vccd1 vccd1 _09622_ sky130_fd_sc_hd__o22a_1
XFILLER_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18721_ _02413_ vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15933_ _08569_ _08577_ vssd1 vssd1 vccd1 vccd1 _08578_ sky130_fd_sc_hd__xnor2_2
X_11056_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _03876_ vssd1 vssd1 vccd1 vccd1 _03878_
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18652_ _02342_ _02347_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _08487_ _08506_ _08508_ vssd1 vssd1 vccd1 vccd1 _08509_ sky130_fd_sc_hd__a21oi_4
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ _10023_ _10025_ vssd1 vssd1 vccd1 vccd1 _10169_ sky130_fd_sc_hd__or2_1
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14815_ _05894_ _07413_ _07516_ _07473_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__a22o_1
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ _02278_ _02279_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__and2b_1
XFILLER_91_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_100 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_100/HI zeros[10]
+ sky130_fd_sc_hd__conb_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _08400_ _08409_ vssd1 vssd1 vccd1 vccd1 _08440_ sky130_fd_sc_hd__xnor2_1
Xtop_ew_algofoogle_111 vssd1 vssd1 vccd1 vccd1 ones[5] top_ew_algofoogle_111/LO sky130_fd_sc_hd__conb_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17534_ _09276_ _08570_ _09417_ _08111_ vssd1 vssd1 vccd1 vccd1 _10100_ sky130_fd_sc_hd__o22a_1
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _05844_ _07477_ _07479_ _07480_ _05800_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__a311o_1
XFILLER_205_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11958_ _04207_ _04708_ _04716_ _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a31o_1
XFILLER_45_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10909_ rbzero.tex_b1\[36\] rbzero.tex_b1\[37\] _03795_ vssd1 vssd1 vccd1 vccd1 _03801_
+ sky130_fd_sc_hd__mux2_1
X_17465_ _10029_ _09902_ _10030_ _10031_ vssd1 vssd1 vccd1 vccd1 _10032_ sky130_fd_sc_hd__a211o_1
XFILLER_205_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14677_ _07407_ _07409_ _07412_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__and3b_1
X_11889_ _04663_ _04665_ _04521_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__a21bo_4
X_19204_ rbzero.spi_registers.new_sky\[5\] rbzero.color_sky\[5\] _02740_ vssd1 vssd1
+ vccd1 vccd1 _02749_ sky130_fd_sc_hd__mux2_1
XFILLER_177_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16416_ _08549_ _08957_ _09060_ vssd1 vssd1 vccd1 vccd1 _09061_ sky130_fd_sc_hd__a21o_2
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13628_ _06360_ _06363_ _06364_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__and3_1
X_17396_ _09961_ _09962_ vssd1 vssd1 vccd1 vccd1 _09963_ sky130_fd_sc_hd__and2_1
XFILLER_38_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19135_ _02702_ vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__clkbuf_1
X_16347_ _08241_ _08247_ vssd1 vssd1 vccd1 vccd1 _08992_ sky130_fd_sc_hd__nor2_1
XFILLER_185_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13559_ _06294_ _06295_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19066_ _02665_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__clkbuf_1
X_16278_ _08867_ _08875_ vssd1 vssd1 vccd1 vccd1 _08923_ sky130_fd_sc_hd__or2_1
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18017_ _08259_ _08157_ _08149_ _08188_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__o22ai_1
XFILLER_173_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15229_ _07821_ _04033_ _07878_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__or3_1
XFILLER_161_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19968_ rbzero.pov.ready_buffer\[41\] _03247_ _03249_ rbzero.debug_overlay.facingX\[-1\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__a221o_1
XFILLER_87_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18919_ _02585_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19899_ _07908_ _03141_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__nor2_1
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20812_ clknet_leaf_66_i_clk _00581_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20743_ clknet_leaf_42_i_clk _00512_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20674_ clknet_leaf_60_i_clk _00458_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_177_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03290_ clknet_0__03290_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03290_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21226_ clknet_leaf_24_i_clk _00995_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21157_ clknet_leaf_68_i_clk _00926_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21088_ net178 _00857_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20039_ _02741_ _03278_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__nor2_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12930_ _05652_ _05659_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nand2_1
XFILLER_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19577__34 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__inv_2
X_12861_ _05481_ _05597_ _05561_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__mux2_2
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _07107_ _07335_ _07336_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__or3b_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _04207_ _04564_ _04572_ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a31o_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _08219_ _08221_ _08224_ vssd1 vssd1 vccd1 vccd1 _08225_ sky130_fd_sc_hd__a21oi_2
XFILLER_14_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ rbzero.wall_tracer.mapY\[5\] _05397_ _05406_ vssd1 vssd1 vccd1 vccd1 _05535_
+ sky130_fd_sc_hd__a21o_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20124__156 clknet_1_1__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__inv_2
XFILLER_42_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _07252_ _07267_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__xnor2_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592__48 clknet_1_0__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__inv_2
X_11743_ _04411_ _04413_ _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__o21a_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _08944_ _08948_ _09826_ vssd1 vssd1 vccd1 vccd1 _09827_ sky130_fd_sc_hd__a21o_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _07162_ _07194_ _07198_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__o21a_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11674_ _04445_ _04449_ _04451_ _04452_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__or4_4
XFILLER_109_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16201_ _08812_ _08844_ vssd1 vssd1 vccd1 vccd1 _08846_ sky130_fd_sc_hd__xor2_1
X_13413_ _06145_ _06149_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__nor2_1
XFILLER_174_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ rbzero.tex_g1\[43\] rbzero.tex_g1\[44\] _03647_ vssd1 vssd1 vccd1 vccd1 _03652_
+ sky130_fd_sc_hd__mux2_1
X_17181_ rbzero.traced_texa\[8\] _09770_ _09771_ rbzero.wall_tracer.visualWallDist\[8\]
+ vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__a22o_1
X_14393_ _06689_ _07072_ _07110_ _07108_ _06675_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__o32ai_1
XFILLER_195_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16132_ _08767_ _08579_ _08727_ _08776_ _08774_ vssd1 vssd1 vccd1 vccd1 _08777_ sky130_fd_sc_hd__o41a_1
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10556_ _03615_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__clkbuf_1
X_13344_ _06078_ _06080_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__or2_1
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16063_ _08704_ _08706_ _08707_ vssd1 vssd1 vccd1 vccd1 _08708_ sky130_fd_sc_hd__a21oi_2
X_10487_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _03569_ vssd1 vssd1 vccd1 vccd1 _03579_
+ sky130_fd_sc_hd__mux2_1
X_13275_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__inv_2
X_15014_ _07678_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__buf_4
X_12226_ _04977_ net16 vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__nand2_1
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12157_ _04907_ _04910_ net68 _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a31o_1
XFILLER_2_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19822_ _03140_ _03143_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__nand2_1
XFILLER_155_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ rbzero.tex_b0\[6\] rbzero.tex_b0\[5\] _03898_ vssd1 vssd1 vccd1 vccd1 _03905_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12088_ net40 _04855_ _04853_ net39 _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__a221o_1
X_16965_ _09587_ _09589_ vssd1 vssd1 vccd1 vccd1 _09605_ sky130_fd_sc_hd__nor2_1
X_19753_ rbzero.pov.spi_buffer\[50\] rbzero.pov.spi_buffer\[51\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03105_ sky130_fd_sc_hd__mux2_1
XFILLER_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15916_ _08482_ _08559_ vssd1 vssd1 vccd1 vccd1 _08561_ sky130_fd_sc_hd__xor2_1
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11039_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _03865_ vssd1 vssd1 vccd1 vccd1 _03869_
+ sky130_fd_sc_hd__mux2_1
X_18704_ _02398_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__buf_4
X_19684_ _03068_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__clkbuf_1
X_16896_ _09520_ _09536_ vssd1 vssd1 vccd1 vccd1 _09537_ sky130_fd_sc_hd__xor2_1
XFILLER_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18635_ _09429_ _09433_ _08356_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a21o_1
XFILLER_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _08129_ _08047_ _08135_ _08491_ vssd1 vssd1 vccd1 vccd1 _08492_ sky130_fd_sc_hd__or4_4
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18566_ _02261_ _02262_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__and2_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15778_ rbzero.wall_tracer.visualWallDist\[5\] _04014_ vssd1 vssd1 vccd1 vccd1 _08423_
+ sky130_fd_sc_hd__nand2_8
XFILLER_45_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17517_ _10080_ _10082_ vssd1 vssd1 vccd1 vccd1 _10083_ sky130_fd_sc_hd__xor2_1
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14729_ _07456_ _07464_ _07459_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__mux2_2
X_18497_ _02084_ _02092_ _02194_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20099__133 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__inv_2
X_17448_ _09955_ _10014_ vssd1 vssd1 vccd1 vccd1 _10015_ sky130_fd_sc_hd__xnor2_2
XFILLER_162_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17379_ _09940_ _09945_ vssd1 vssd1 vccd1 vccd1 _09946_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19118_ _02693_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19049_ _02656_ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21011_ clknet_leaf_12_i_clk _00780_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20726_ clknet_leaf_83_i_clk _00495_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20657_ clknet_leaf_56_i_clk _00441_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10410_ _03536_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _04160_ gpout0.hpos\[5\] _04022_ _04161_ _04169_ vssd1 vssd1 vccd1 vccd1
+ _04170_ sky130_fd_sc_hd__o221a_1
X_20588_ _07683_ _07692_ _07691_ _07831_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__a31o_1
XFILLER_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10341_ _03500_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13060_ _05795_ _05796_ _05743_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__a21o_1
XFILLER_155_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12011_ _04210_ _04781_ _04785_ _04371_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a211o_1
X_21209_ clknet_leaf_26_i_clk _00978_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16750_ _09391_ _08356_ _09389_ vssd1 vssd1 vccd1 vccd1 _09392_ sky130_fd_sc_hd__o21ai_1
X_13962_ _06698_ _06690_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__nor2_2
XFILLER_4_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15701_ _08076_ _08085_ _08106_ vssd1 vssd1 vccd1 vccd1 _08346_ sky130_fd_sc_hd__o21ba_1
X_12913_ _05601_ _05606_ _05638_ _05649_ _05628_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__o41a_2
XFILLER_111_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16681_ _09321_ _09323_ vssd1 vssd1 vccd1 vccd1 _09324_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13893_ _06579_ _06628_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__nand2_1
XFILLER_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18420_ _01807_ _01810_ _01927_ _01925_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__a31oi_1
X_15632_ _08276_ _08008_ vssd1 vssd1 vccd1 vccd1 _08277_ sky130_fd_sc_hd__nor2_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12844_ rbzero.wall_tracer.visualWallDist\[-5\] _05570_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05581_ sky130_fd_sc_hd__a21o_1
XFILLER_74_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18351_ _01988_ _01989_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__nand2_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _07560_ _07562_ _07564_ _08171_ vssd1 vssd1 vccd1 vccd1 _08208_ sky130_fd_sc_hd__nor4_2
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _05511_ _05515_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__or2_1
XFILLER_199_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.stepDistX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _09873_ sky130_fd_sc_hd__nand2_1
XFILLER_202_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _07245_ _07244_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__and2b_1
X_18282_ _01737_ _09693_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__nor2_1
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ rbzero.debug_overlay.playerY\[5\] _04444_ _04439_ _04465_ rbzero.debug_overlay.playerY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__a32o_1
X_15494_ _08109_ _08042_ vssd1 vssd1 vccd1 vccd1 _08139_ sky130_fd_sc_hd__or2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17233_ _05243_ _09781_ _09811_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14445_ _07175_ _07180_ _07181_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__o21a_1
X_11657_ _04415_ _04430_ _04417_ _04022_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__or4b_2
XFILLER_35_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10608_ _03642_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__clkbuf_1
X_17164_ rbzero.traced_texa\[-6\] _09768_ _09767_ rbzero.wall_tracer.visualWallDist\[-6\]
+ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__a22o_1
XFILLER_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ _06689_ _06760_ _07110_ _07108_ _06675_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__o32a_1
X_11588_ rbzero.tex_r1\[29\] rbzero.tex_r1\[28\] _04342_ vssd1 vssd1 vccd1 vccd1 _04367_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16115_ _08756_ _08758_ _08759_ vssd1 vssd1 vccd1 vccd1 _08760_ sky130_fd_sc_hd__a21oi_2
XFILLER_156_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13327_ _06058_ _06062_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10539_ _03606_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__clkbuf_1
X_17095_ _09605_ _09606_ _09734_ vssd1 vssd1 vccd1 vccd1 _09735_ sky130_fd_sc_hd__nor3_1
XFILLER_182_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16046_ _08662_ _08690_ vssd1 vssd1 vccd1 vccd1 _08691_ sky130_fd_sc_hd__nand2_1
XFILLER_131_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13258_ _05994_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__buf_2
XFILLER_142_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12209_ _04323_ _04962_ _04978_ net68 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__a22o_1
XFILLER_170_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _05807_ _05858_ _05871_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19805_ _03131_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17997_ _01615_ _01630_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__nor2_1
X_20399__24 clknet_1_0__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__inv_2
XFILLER_85_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03305_ clknet_0__03305_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03305_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16948_ _09347_ _09450_ _09588_ vssd1 vssd1 vccd1 vccd1 _09589_ sky130_fd_sc_hd__a21oi_1
X_19736_ rbzero.pov.spi_buffer\[42\] rbzero.pov.spi_buffer\[43\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03096_ sky130_fd_sc_hd__mux2_1
XFILLER_38_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16879_ _09407_ _09414_ _09519_ vssd1 vssd1 vccd1 vccd1 _09520_ sky130_fd_sc_hd__a21o_1
X_19667_ rbzero.pov.spi_buffer\[9\] rbzero.pov.spi_buffer\[10\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03060_ sky130_fd_sc_hd__mux2_1
XFILLER_42_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18618_ _02312_ _02314_ _05204_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a21o_1
XFILLER_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20107__140 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__inv_2
XFILLER_206_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18549_ _02241_ _02245_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__xor2_1
XFILLER_205_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21560_ net481 _01329_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20511_ rbzero.traced_texa\[4\] rbzero.texV\[4\] vssd1 vssd1 vccd1 vccd1 _03407_
+ sky130_fd_sc_hd__nor2_1
X_21491_ net412 _01260_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20442_ _03343_ _03345_ _03344_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__o21bai_1
XFILLER_118_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20153__182 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__inv_2
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10890_ rbzero.tex_b1\[45\] rbzero.tex_b1\[46\] _03784_ vssd1 vssd1 vccd1 vccd1 _03791_
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12560_ _05313_ _05287_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__nor2_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11511_ _04290_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__clkbuf_8
XFILLER_197_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20709_ clknet_leaf_71_i_clk _00000_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12491_ rbzero.wall_tracer.trackDistY\[-9\] _05240_ rbzero.wall_tracer.trackDistY\[-10\]
+ _05241_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__o221a_1
XFILLER_156_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14230_ _06888_ _06966_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__nand2_1
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11442_ _04136_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20236__257 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__inv_2
XFILLER_153_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11373_ rbzero.row_render.size\[7\] _04152_ rbzero.row_render.size\[8\] vssd1 vssd1
+ vccd1 vccd1 _04153_ sky130_fd_sc_hd__o21a_1
XFILLER_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14161_ _06894_ _06896_ _06897_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10324_ _03491_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__clkbuf_1
X_13112_ _05718_ _05734_ _05803_ _05721_ _05777_ _05801_ vssd1 vssd1 vccd1 vccd1 _05849_
+ sky130_fd_sc_hd__mux4_1
XFILLER_180_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14092_ _06804_ _06828_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17920_ _08802_ _09693_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__nor2_1
XFILLER_140_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _05695_ _05702_ _05677_ _05762_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__or4_1
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17851_ rbzero.wall_tracer.trackDistX\[3\] rbzero.wall_tracer.stepDistX\[3\] vssd1
+ vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__or2_1
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16802_ _09442_ _09443_ vssd1 vssd1 vccd1 vccd1 _09444_ sky130_fd_sc_hd__xor2_1
XFILLER_182_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17782_ _10215_ _10224_ _10222_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14994_ _07667_ vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16733_ _09372_ _09374_ vssd1 vssd1 vccd1 vccd1 _09375_ sky130_fd_sc_hd__nor2_1
XFILLER_47_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19521_ _03913_ _02997_ _02998_ _07695_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a31o_1
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _06675_ _06668_ _06681_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__o21ba_1
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19452_ _07831_ _02925_ _02926_ _02934_ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__o31ai_1
X_16664_ _09145_ _09147_ vssd1 vssd1 vccd1 vccd1 _09307_ sky130_fd_sc_hd__nor2_1
X_13876_ _06560_ _06601_ _06603_ _06612_ vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__a211oi_2
XFILLER_62_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18403_ _02060_ _02101_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__xnor2_2
X_15615_ _08259_ _08226_ _08244_ vssd1 vssd1 vccd1 vccd1 _08260_ sky130_fd_sc_hd__or3_1
X_19383_ _02868_ _02869_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nand2_1
X_12827_ _03953_ _04030_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__nor2_1
X_16595_ _09210_ _09237_ vssd1 vssd1 vccd1 vccd1 _09238_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18334_ _02031_ _02032_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__nor2_1
X_15546_ _08177_ _07989_ vssd1 vssd1 vccd1 vccd1 _08191_ sky130_fd_sc_hd__nor2_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ rbzero.map_rom.f2 _05496_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__nor2_1
XFILLER_203_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18265_ _01932_ _01964_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__xor2_1
X_11709_ rbzero.debug_overlay.facingY\[10\] _04453_ _04487_ vssd1 vssd1 vccd1 vccd1
+ _04488_ sky130_fd_sc_hd__a21oi_1
X_15477_ _08120_ _08121_ vssd1 vssd1 vccd1 vccd1 _08122_ sky130_fd_sc_hd__nand2_1
X_12689_ _05420_ _05431_ _05419_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__a21o_1
X_17216_ rbzero.wall_tracer.mapX\[10\] _05525_ vssd1 vssd1 vccd1 vccd1 _09797_ sky130_fd_sc_hd__xor2_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ _06067_ _06668_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__or2_1
X_18196_ _01817_ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ rbzero.row_render.size\[9\] _09762_ _07560_ _07756_ vssd1 vssd1 vccd1 vccd1
+ _00537_ sky130_fd_sc_hd__a22o_1
X_14359_ _07031_ _07033_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__nor2_1
XFILLER_143_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17078_ _09692_ _09717_ vssd1 vssd1 vccd1 vccd1 _09718_ sky130_fd_sc_hd__xnor2_4
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16029_ _08019_ vssd1 vssd1 vccd1 vccd1 _08674_ sky130_fd_sc_hd__clkbuf_4
XFILLER_115_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19719_ rbzero.pov.spi_buffer\[34\] rbzero.pov.spi_buffer\[35\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03087_ sky130_fd_sc_hd__mux2_1
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20991_ clknet_leaf_14_i_clk _00760_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03319_ _03319_ vssd1 vssd1 vccd1 vccd1 clknet_0__03319_ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21612_ net129 _01381_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21543_ net464 _01312_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21474_ net395 _01243_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[53\] sky130_fd_sc_hd__dfxtp_1
X_20425_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 _03335_
+ sky130_fd_sc_hd__nand2_1
XFILLER_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03041_ clknet_0__03041_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03041_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11991_ rbzero.tex_b1\[3\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__and3_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ _06440_ _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__xor2_1
X_10942_ _03818_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13661_ _06365_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__or2_1
XFILLER_95_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10873_ rbzero.tex_b1\[53\] rbzero.tex_b1\[54\] _03773_ vssd1 vssd1 vccd1 vccd1 _03782_
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15400_ _07945_ _08044_ vssd1 vssd1 vccd1 vccd1 _08045_ sky130_fd_sc_hd__or2_1
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _05308_ _05312_ _05318_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__o21a_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _09022_ _09024_ vssd1 vssd1 vccd1 vccd1 _09025_ sky130_fd_sc_hd__xor2_4
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _06303_ _06328_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__xnor2_1
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15331_ _07925_ _07974_ _07975_ _05207_ vssd1 vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__a211o_2
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12543_ rbzero.debug_overlay.facingY\[-3\] rbzero.wall_tracer.rayAddendY\[5\] vssd1
+ vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__nand2_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18050_ _01736_ _01751_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15262_ rbzero.debug_overlay.playerY\[-6\] _07905_ vssd1 vssd1 vccd1 vccd1 _07907_
+ sky130_fd_sc_hd__nand2_1
X_12474_ _05219_ _05227_ _05228_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__o21a_1
Xclkbuf_1_0__f__03308_ clknet_0__03308_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03308_
+ sky130_fd_sc_hd__clkbuf_16
X_17001_ _09245_ _08159_ vssd1 vssd1 vccd1 vccd1 _09641_ sky130_fd_sc_hd__nor2_1
X_14213_ _06666_ _06690_ _06921_ _06919_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__o31a_1
XFILLER_184_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ rbzero.floor_leak\[5\] _04116_ _04133_ _04134_ _04204_ vssd1 vssd1 vccd1
+ vccd1 _04205_ sky130_fd_sc_hd__a221o_1
X_15193_ _07843_ _07844_ _07841_ _07842_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__a211o_1
XANTENNA_7 _07524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ _06856_ _06879_ _06880_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__a21oi_2
XFILLER_4_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ _04127_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__clkbuf_4
XFILLER_126_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10307_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__clkbuf_4
X_14075_ _06803_ _06810_ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__nor2_1
X_18952_ rbzero.pov.spi_buffer\[9\] rbzero.pov.ready_buffer\[9\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02606_ sky130_fd_sc_hd__mux2_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11287_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] vssd1 vssd1
+ vccd1 vccd1 _04067_ sky130_fd_sc_hd__nand2_1
XFILLER_112_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17903_ _01604_ _01605_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__nor2_1
X_13026_ _05761_ _05762_ _05748_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__and3_1
XFILLER_6_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18883_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_cmd\[2\]
+ rbzero.spi_registers.spi_cmd\[0\] vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__and4bb_1
XFILLER_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17834_ _01535_ _01537_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__xor2_1
XFILLER_117_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17765_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__and2_1
XFILLER_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14977_ _00008_ _07536_ _07658_ vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19504_ rbzero.debug_overlay.vplaneY\[-1\] _02961_ vssd1 vssd1 vccd1 vccd1 _02983_
+ sky130_fd_sc_hd__nand2_1
X_16716_ _09356_ _09357_ vssd1 vssd1 vccd1 vccd1 _09358_ sky130_fd_sc_hd__xnor2_1
X_13928_ _06659_ _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__nand2_1
XFILLER_207_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17696_ _10110_ _09973_ vssd1 vssd1 vccd1 vccd1 _10261_ sky130_fd_sc_hd__nor2_1
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16647_ _08215_ _08519_ _08985_ _09138_ vssd1 vssd1 vccd1 vccd1 _09290_ sky130_fd_sc_hd__or4_1
XFILLER_23_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19435_ _02908_ _02909_ _02918_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__o21ai_1
X_13859_ _06564_ _06594_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__or2_1
XFILLER_179_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16578_ _09161_ _09219_ vssd1 vssd1 vccd1 vccd1 _09221_ sky130_fd_sc_hd__or2_1
X_19366_ _02854_ _02842_ _02841_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_65_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18317_ rbzero.wall_tracer.trackDistX\[7\] rbzero.wall_tracer.stepDistX\[7\] vssd1
+ vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__or2_1
XFILLER_37_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15529_ _07894_ _05342_ _08173_ _07970_ vssd1 vssd1 vccd1 vccd1 _08174_ sky130_fd_sc_hd__o211a_1
XFILLER_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19297_ _02804_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__clkbuf_1
X_18248_ _01946_ _01947_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__and2_1
XFILLER_176_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20219__241 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__inv_2
XFILLER_198_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18179_ _10110_ _10266_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__nor2_1
XFILLER_128_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21190_ clknet_leaf_22_i_clk _00959_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20072_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__buf_1
XFILLER_106_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_18_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20265__283 clknet_1_1__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__inv_2
XFILLER_39_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20974_ clknet_leaf_12_i_clk _00743_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21526_ net447 _01295_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21457_ net378 _01226_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11210_ _03970_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__and2_1
X_12190_ net15 vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__buf_2
X_20408_ gpout5.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__nor2_1
XFILLER_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21388_ net309 _01157_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ rbzero.debug_overlay.playerY\[0\] vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__inv_2
XFILLER_150_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput55 net55 vssd1 vssd1 vccd1 vccd1 o_gpout[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_122_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput66 net66 vssd1 vssd1 vccd1 vccd1 o_rgb[7] sky130_fd_sc_hd__buf_2
XFILLER_153_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11072_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _03876_ vssd1 vssd1 vccd1 vccd1 _03886_
+ sky130_fd_sc_hd__mux2_1
XFILLER_163_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14900_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.trackDistX\[-7\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__mux2_1
X_20348__358 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__inv_2
XFILLER_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15880_ _08522_ _08523_ _08524_ vssd1 vssd1 vccd1 vccd1 _08525_ sky130_fd_sc_hd__o21ba_1
XFILLER_49_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ rbzero.wall_tracer.stepDistY\[0\] _07461_ vssd1 vssd1 vccd1 vccd1 _07556_
+ sky130_fd_sc_hd__nor2_1
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ _09980_ _10115_ vssd1 vssd1 vccd1 vccd1 _10116_ sky130_fd_sc_hd__xnor2_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14762_ _05884_ _07492_ _07495_ vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__a21o_1
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ rbzero.tex_b1\[29\] rbzero.tex_b1\[28\] _04342_ vssd1 vssd1 vccd1 vccd1 _04749_
+ sky130_fd_sc_hd__mux2_1
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16501_ _09132_ _09144_ vssd1 vssd1 vccd1 vccd1 _09145_ sky130_fd_sc_hd__xnor2_2
XFILLER_189_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13713_ _06041_ _06449_ _06407_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__mux2_1
XFILLER_44_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17481_ _10045_ _10046_ vssd1 vssd1 vccd1 vccd1 _10047_ sky130_fd_sc_hd__nor2_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _03809_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14693_ _05779_ _07428_ _07429_ _05892_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__o211a_1
X_19220_ _02759_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__clkbuf_1
X_16432_ _09074_ _09075_ _09076_ vssd1 vssd1 vccd1 vccd1 _09077_ sky130_fd_sc_hd__a21o_1
XFILLER_177_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13644_ _05988_ _06380_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__xnor2_1
X_10856_ _03646_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19151_ rbzero.spi_registers.new_other\[8\] _02712_ vssd1 vssd1 vccd1 vccd1 _02716_
+ sky130_fd_sc_hd__or2_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16363_ _09006_ _09007_ vssd1 vssd1 vccd1 vccd1 _09008_ sky130_fd_sc_hd__and2_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13575_ _05823_ _05961_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__or2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ rbzero.tex_g0\[31\] rbzero.tex_g0\[30\] _03729_ vssd1 vssd1 vccd1 vccd1 _03737_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18102_ _01784_ _01686_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__or2b_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _07958_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__buf_4
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19082_ _02673_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__clkbuf_1
X_12526_ _03912_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__nor2_1
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16294_ _08803_ _08804_ _08807_ _08938_ vssd1 vssd1 vccd1 vccd1 _08939_ sky130_fd_sc_hd__a211oi_1
XFILLER_121_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18033_ _01622_ _01629_ _01734_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__a21o_1
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20093__128 clknet_1_0__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__inv_2
X_15245_ _04035_ _07891_ vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__and2_1
X_12457_ rbzero.wall_tracer.trackDistX\[11\] vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__inv_2
XFILLER_126_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11408_ rbzero.row_render.size\[3\] _04149_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__nand2_1
X_15176_ _04033_ _04027_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__nand2_8
X_12388_ net40 _05145_ _05143_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__and3_1
XFILLER_153_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ _06769_ _06667_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__nor2_1
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11339_ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__clkbuf_4
XFILLER_4_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19984_ rbzero.pov.ready_buffer\[11\] _03246_ _03248_ rbzero.debug_overlay.vplaneX\[-9\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__a221o_1
X_14058_ _06789_ _06793_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__or2b_1
X_18935_ rbzero.pov.spi_buffer\[1\] rbzero.pov.ready_buffer\[1\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02597_ sky130_fd_sc_hd__mux2_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13009_ _05690_ _05702_ _05683_ _05745_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__or4_1
XFILLER_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18866_ _02537_ _02538_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17817_ _01519_ _01520_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__xnor2_1
XFILLER_94_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18797_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.stepDistY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__nor2_1
XFILLER_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17748_ _01443_ _01444_ _01450_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__and3_1
XFILLER_78_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17679_ _08802_ _09552_ vssd1 vssd1 vccd1 vccd1 _10244_ sky130_fd_sc_hd__nor2_2
XFILLER_165_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19418_ rbzero.wall_tracer.rayAddendY\[1\] _07695_ _02902_ _07703_ vssd1 vssd1 vccd1
+ vccd1 _02903_ sky130_fd_sc_hd__a22o_1
XFILLER_168_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20690_ clknet_leaf_55_i_clk _00474_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19349_ _07728_ _02838_ _02839_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__a21o_1
XFILLER_149_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21311_ net232 _01080_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21242_ clknet_leaf_91_i_clk _01011_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21173_ clknet_leaf_78_i_clk _00942_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20957_ clknet_leaf_94_i_clk _00726_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _03696_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__clkbuf_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11690_ rbzero.debug_overlay.vplaneX\[-9\] _04458_ _04461_ _04468_ vssd1 vssd1 vccd1
+ vccd1 _04469_ sky130_fd_sc_hd__a211o_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20888_ clknet_leaf_86_i_clk _00657_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_186_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ _03660_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13360_ _06094_ _06095_ _06096_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__nand3_1
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10572_ _03623_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12311_ net24 net25 net66 _05068_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__or4_1
X_21509_ net430 _01278_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13291_ _05855_ _06010_ _06025_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__a22o_1
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15030_ _04028_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__buf_4
X_12242_ _04867_ _04964_ net47 vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ _04154_ _03477_ net8 vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__mux2_1
XFILLER_162_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11124_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__buf_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16981_ _05211_ _09350_ vssd1 vssd1 vccd1 vccd1 _09621_ sky130_fd_sc_hd__nor2_1
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18720_ rbzero.wall_tracer.trackDistY\[-10\] _02412_ _02399_ vssd1 vssd1 vccd1 vccd1
+ _02413_ sky130_fd_sc_hd__mux2_1
XFILLER_95_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15932_ _08570_ _08128_ _08571_ _08576_ vssd1 vssd1 vccd1 vccd1 _08577_ sky130_fd_sc_hd__o31a_1
XFILLER_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11055_ _03877_ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_27_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18651_ _02345_ _02346_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__xnor2_1
X_15863_ _08154_ _08507_ vssd1 vssd1 vccd1 vccd1 _08508_ sky130_fd_sc_hd__nand2_1
XFILLER_49_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ _10023_ _10025_ vssd1 vssd1 vccd1 vccd1 _10168_ sky130_fd_sc_hd__and2_1
X_14814_ _07542_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__clkbuf_1
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18582_ _02272_ _02277_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__or2_1
X_15794_ _08412_ _08438_ vssd1 vssd1 vccd1 vccd1 _08439_ sky130_fd_sc_hd__xnor2_2
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_101 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_101/HI zeros[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_188_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_112 vssd1 vssd1 vccd1 vccd1 ones[6] top_ew_algofoogle_112/LO sky130_fd_sc_hd__conb_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ _09668_ _09417_ vssd1 vssd1 vccd1 vccd1 _10099_ sky130_fd_sc_hd__nor2_2
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14745_ _07384_ _07401_ _05844_ _05952_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__o211a_1
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _04244_ _04724_ _04732_ _04116_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a31o_1
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10908_ _03800_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__clkbuf_1
X_17464_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] vssd1
+ vssd1 vccd1 vccd1 _10031_ sky130_fd_sc_hd__and2_1
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14676_ _07407_ _07410_ _07412_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__o21ba_2
XFILLER_189_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11888_ _04206_ _04664_ _04314_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16415_ _09059_ _08547_ vssd1 vssd1 vccd1 vccd1 _09060_ sky130_fd_sc_hd__xnor2_2
X_19203_ rbzero.color_sky\[4\] _02740_ _02748_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__a21o_1
X_13627_ _06078_ _05982_ _06361_ _06362_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__o211ai_1
X_17395_ _09661_ _08356_ _09960_ vssd1 vssd1 vccd1 vccd1 _09962_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10839_ _03764_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__clkbuf_1
X_20101__135 clknet_1_1__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__inv_2
XFILLER_34_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16346_ _08976_ _08990_ vssd1 vssd1 vccd1 vccd1 _08991_ sky130_fd_sc_hd__xnor2_2
X_19134_ rbzero.spi_registers.sclk_buffer\[1\] rbzero.spi_registers.sclk_buffer\[2\]
+ _02695_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__mux2_1
X_13558_ _05888_ _05923_ _06116_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__and3_1
XFILLER_34_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19065_ rbzero.pov.spi_buffer\[63\] rbzero.pov.ready_buffer\[63\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02665_ sky130_fd_sc_hd__mux2_1
X_12509_ rbzero.wall_tracer.trackDistX\[3\] vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__inv_2
X_16277_ _08912_ _08913_ _08920_ _08921_ vssd1 vssd1 vccd1 vccd1 _08922_ sky130_fd_sc_hd__and4b_1
XFILLER_195_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13489_ _06197_ _06198_ _06224_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__or3_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18016_ _08259_ _08188_ _08157_ _08149_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__or4_1
X_15228_ _07730_ _07854_ vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__nor2_1
XFILLER_133_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15159_ _07803_ _07808_ _07813_ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__o21a_1
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19967_ rbzero.pov.ready_buffer\[40\] _03240_ _03243_ rbzero.debug_overlay.facingX\[-2\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__o221a_1
XFILLER_45_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18918_ _02583_ _02584_ _02574_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__and3b_1
XFILLER_45_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19898_ rbzero.debug_overlay.playerY\[-7\] _03198_ _03202_ _03157_ vssd1 vssd1 vccd1
+ vccd1 _00991_ sky130_fd_sc_hd__o211a_1
XFILLER_80_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18849_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.stepDistY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__nand2_1
XFILLER_83_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20811_ clknet_leaf_66_i_clk _00580_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20742_ clknet_leaf_42_i_clk _00511_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20673_ clknet_leaf_48_i_clk _00457_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[2\]
+ sky130_fd_sc_hd__dfxtp_4
X_20377__384 clknet_1_0__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__inv_2
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20076__112 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__inv_2
XFILLER_177_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21225_ clknet_leaf_24_i_clk _00994_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_176_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21156_ clknet_leaf_85_i_clk _00925_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21087_ net177 _00856_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20038_ _04990_ _04989_ _04037_ _02705_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__and4_1
XFILLER_19_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ rbzero.wall_tracer.visualWallDist\[-8\] _05353_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__mux2_1
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _04121_ _04580_ _04588_ _04116_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__a31o_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12791_ rbzero.wall_tracer.mapY\[6\] _05397_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__xor2_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14530_ _07259_ _07266_ _07264_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__a21oi_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _04519_ _04520_ _04021_ _04323_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__a211oi_4
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _07195_ _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__or2b_1
XFILLER_202_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _04432_ _04448_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__nor2_1
XFILLER_168_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16200_ _08812_ _08844_ vssd1 vssd1 vccd1 vccd1 _08845_ sky130_fd_sc_hd__or2_1
XFILLER_70_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13412_ _06147_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__and2b_1
X_10624_ _03651_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__clkbuf_1
X_17180_ _07679_ vssd1 vssd1 vccd1 vccd1 _09771_ sky130_fd_sc_hd__clkbuf_4
X_14392_ _07111_ _07128_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__or2_1
XFILLER_183_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _08774_ _08775_ vssd1 vssd1 vccd1 vccd1 _08776_ sky130_fd_sc_hd__nand2_1
XFILLER_127_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13343_ _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__clkbuf_4
XFILLER_194_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10555_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _03613_ vssd1 vssd1 vccd1 vccd1 _03615_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16062_ _08702_ _08703_ vssd1 vssd1 vccd1 vccd1 _08707_ sky130_fd_sc_hd__and2_1
X_13274_ _05946_ _05877_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10486_ _03578_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15013_ _07676_ _07677_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__nor2_1
X_12225_ _04986_ _04994_ net19 vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__and3b_1
XFILLER_185_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19821_ _03138_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__clkbuf_4
X_12156_ net46 _04918_ _04922_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a22o_1
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03321_ clknet_0__03321_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03321_
+ sky130_fd_sc_hd__clkbuf_16
X_11107_ _03904_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__clkbuf_1
X_19752_ _03104_ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12087_ net38 _04857_ _04838_ net48 vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__a22o_1
X_16964_ rbzero.wall_tracer.texu\[4\] _09085_ _04035_ _09604_ vssd1 vssd1 vccd1 vccd1
+ _00515_ sky130_fd_sc_hd__o211a_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18703_ _05203_ _09283_ _05282_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__o21a_2
X_15915_ _07959_ _08042_ vssd1 vssd1 vccd1 vccd1 _08560_ sky130_fd_sc_hd__nor2_1
X_11038_ _03868_ vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__clkbuf_1
X_19683_ rbzero.pov.spi_buffer\[17\] rbzero.pov.spi_buffer\[18\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03068_ sky130_fd_sc_hd__mux2_1
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16895_ _09528_ _09535_ vssd1 vssd1 vccd1 vccd1 _09536_ sky130_fd_sc_hd__xnor2_2
X_18634_ _02326_ _02329_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _08124_ _08490_ vssd1 vssd1 vccd1 vccd1 _08491_ sky130_fd_sc_hd__and2_4
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18565_ _01739_ _09027_ _02260_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__o21ai_1
XFILLER_75_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15777_ _08416_ _08420_ _08421_ vssd1 vssd1 vccd1 vccd1 _08422_ sky130_fd_sc_hd__a21o_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12989_ _05657_ _05658_ _05663_ _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__or4b_1
XFILLER_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17516_ _09939_ _09946_ _10081_ vssd1 vssd1 vccd1 vccd1 _10082_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14728_ _07463_ _07424_ _07433_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__mux2_1
X_18496_ _02085_ _01985_ _02091_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__a21oi_1
XFILLER_162_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17447_ _10011_ _10013_ vssd1 vssd1 vccd1 vccd1 _10014_ sky130_fd_sc_hd__xnor2_1
X_14659_ _07103_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__clkinv_2
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17378_ _09943_ _09944_ vssd1 vssd1 vccd1 vccd1 _09945_ sky130_fd_sc_hd__xor2_1
XFILLER_203_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19117_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[2\] _02690_
+ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__mux2_1
X_16329_ _08972_ _08973_ vssd1 vssd1 vccd1 vccd1 _08974_ sky130_fd_sc_hd__or2b_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19048_ rbzero.pov.spi_buffer\[55\] rbzero.pov.ready_buffer\[55\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02656_ sky130_fd_sc_hd__mux2_1
XFILLER_106_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21010_ clknet_leaf_12_i_clk _00779_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20725_ clknet_leaf_83_i_clk _00494_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20656_ clknet_leaf_52_i_clk _00440_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20587_ _07683_ _07692_ _07691_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__a21oi_1
X_10340_ rbzero.tex_r1\[48\] rbzero.tex_r1\[49\] _03494_ vssd1 vssd1 vccd1 vccd1 _03500_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _04782_ _04783_ _04784_ _04266_ _04229_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__o221a_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21208_ clknet_leaf_29_i_clk _00977_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21139_ clknet_leaf_97_i_clk _00908_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20130__161 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__inv_2
XFILLER_171_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13961_ _06134_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__clkbuf_4
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15700_ _08343_ _08344_ vssd1 vssd1 vccd1 vccd1 _08345_ sky130_fd_sc_hd__or2_1
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12912_ _05640_ _05642_ _05645_ _05648_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__or4_2
X_16680_ _09160_ _09180_ _09322_ vssd1 vssd1 vccd1 vccd1 _09323_ sky130_fd_sc_hd__a21boi_1
XFILLER_47_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13892_ _06579_ _06628_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__or2_1
XFILLER_59_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12843_ rbzero.wall_tracer.rcp_sel\[2\] _05347_ _05348_ vssd1 vssd1 vccd1 vccd1 _05580_
+ sky130_fd_sc_hd__and3_1
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _08269_ _08275_ _07990_ vssd1 vssd1 vccd1 vccd1 _08276_ sky130_fd_sc_hd__mux2_2
XFILLER_34_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18350_ _02047_ _02048_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15562_ rbzero.wall_tracer.stepDistY\[3\] vssd1 vssd1 vccd1 vccd1 _08207_ sky130_fd_sc_hd__inv_2
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ rbzero.map_rom.i_col\[4\] _05512_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__xor2_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _07233_ _07249_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__xnor2_1
X_17301_ rbzero.wall_tracer.trackDistX\[-4\] rbzero.wall_tracer.stepDistX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _09872_ sky130_fd_sc_hd__nor2_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ rbzero.debug_overlay.playerY\[-3\] _04463_ _04502_ _04503_ vssd1 vssd1 vccd1
+ vccd1 _04504_ sky130_fd_sc_hd__a211o_1
XFILLER_202_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18281_ _01756_ _01881_ _01980_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a21o_1
X_15493_ _08115_ _08116_ vssd1 vssd1 vccd1 vccd1 _08138_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14444_ _07172_ _07174_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__nand2_1
X_17232_ _05413_ _09808_ _09810_ vssd1 vssd1 vccd1 vccd1 _09811_ sky130_fd_sc_hd__and3_1
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11656_ _04420_ _04428_ _04433_ _04434_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__or4_1
XFILLER_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10607_ rbzero.tex_g1\[51\] rbzero.tex_g1\[52\] _03635_ vssd1 vssd1 vccd1 vccd1 _03642_
+ sky130_fd_sc_hd__mux2_1
X_17163_ rbzero.traced_texa\[-7\] _09768_ _09767_ rbzero.wall_tracer.visualWallDist\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__a22o_1
XFILLER_7_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14375_ _07110_ _07111_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__xor2_1
X_11587_ _04364_ _04365_ _04329_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__mux2_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16114_ _08740_ _08755_ vssd1 vssd1 vccd1 vccd1 _08759_ sky130_fd_sc_hd__nor2_1
XFILLER_127_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13326_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__inv_2
XFILLER_183_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10538_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _03602_ vssd1 vssd1 vccd1 vccd1 _03606_
+ sky130_fd_sc_hd__mux2_1
X_17094_ _09474_ _09733_ vssd1 vssd1 vccd1 vccd1 _09734_ sky130_fd_sc_hd__xor2_1
XFILLER_7_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16045_ _08659_ _08661_ vssd1 vssd1 vccd1 vccd1 _08690_ sky130_fd_sc_hd__or2_1
X_13257_ _05979_ _05909_ _05900_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__or3b_1
X_10469_ rbzero.tex_r0\[54\] rbzero.tex_r0\[53\] _03569_ vssd1 vssd1 vccd1 vccd1 _03570_
+ sky130_fd_sc_hd__mux2_1
XFILLER_170_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20213__236 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__inv_2
XFILLER_142_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12208_ net15 net14 vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__and2b_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13188_ _05807_ _05924_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__nand2_1
XFILLER_151_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19804_ net50 rbzero.pov.ss_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__mux2_1
X_12139_ net8 vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__clkbuf_4
XFILLER_96_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17996_ _01591_ _01606_ _01604_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a21o_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03304_ clknet_0__03304_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03304_
+ sky130_fd_sc_hd__clkbuf_16
X_19735_ _03095_ vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16947_ _09448_ _09449_ vssd1 vssd1 vccd1 vccd1 _09588_ sky130_fd_sc_hd__nor2_1
XFILLER_93_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19666_ _03047_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__clkbuf_4
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16878_ _09408_ _09413_ vssd1 vssd1 vccd1 vccd1 _09519_ sky130_fd_sc_hd__and2b_1
XFILLER_77_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18617_ _02125_ _02128_ _02222_ _02223_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__a31o_1
X_15829_ _08008_ _07941_ vssd1 vssd1 vccd1 vccd1 _08474_ sky130_fd_sc_hd__nor2_1
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18548_ _02242_ _02244_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18479_ _01939_ _02071_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__nand2_1
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20510_ _03401_ _03403_ _03402_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__a21boi_1
X_21490_ net411 _01259_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20441_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] vssd1 vssd1 vccd1 vccd1 _03348_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19619__72 clknet_1_0__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__inv_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20188__213 clknet_1_0__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__inv_2
XFILLER_130_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19634__86 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__inv_2
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11510_ _04129_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__clkbuf_8
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20708_ clknet_leaf_47_i_clk _00015_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12490_ rbzero.wall_tracer.trackDistY\[-10\] _05241_ rbzero.wall_tracer.trackDistY\[-11\]
+ _05242_ _05244_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__a221o_1
XFILLER_106_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11441_ _04135_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__clkbuf_4
X_20639_ clknet_leaf_63_i_clk _00423_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14160_ _06864_ _06895_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__and2_1
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11372_ rbzero.row_render.size\[6\] _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__and2_1
XFILLER_192_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ _05838_ _05843_ _05820_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__mux2_1
X_10323_ rbzero.tex_r1\[56\] rbzero.tex_r1\[57\] _03483_ vssd1 vssd1 vccd1 vccd1 _03491_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14091_ _06776_ _06662_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__nor2_1
XFILLER_4_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13042_ _05778_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__buf_2
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17850_ rbzero.wall_tracer.trackDistX\[3\] rbzero.wall_tracer.stepDistX\[3\] vssd1
+ vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__nand2_1
XFILLER_26_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16801_ _09303_ _09305_ vssd1 vssd1 vccd1 vccd1 _09443_ sky130_fd_sc_hd__and2_1
XFILLER_121_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17781_ _01472_ _01484_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__xnor2_1
X_14993_ rbzero.wall_tracer.stepDistX\[3\] _07564_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07667_ sky130_fd_sc_hd__mux2_1
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19520_ _02983_ _02987_ _02996_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__a21o_1
X_16732_ _09223_ _09230_ _09373_ vssd1 vssd1 vccd1 vccd1 _09374_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13944_ _06680_ _06677_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__nor2_1
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19451_ rbzero.wall_tracer.rayAddendY\[3\] _07855_ _02932_ _02933_ vssd1 vssd1 vccd1
+ vccd1 _02934_ sky130_fd_sc_hd__a22oi_1
X_16663_ _09303_ _09304_ _09275_ vssd1 vssd1 vccd1 vccd1 _09306_ sky130_fd_sc_hd__a21o_1
XFILLER_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13875_ _06605_ _06611_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__nor2_4
X_18402_ _02062_ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__xnor2_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12826_ _05562_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__buf_2
X_15614_ _08175_ _08176_ vssd1 vssd1 vccd1 vccd1 _08259_ sky130_fd_sc_hd__nand2_4
X_19382_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__nand2_1
X_16594_ _09222_ _09236_ vssd1 vssd1 vccd1 vccd1 _09237_ sky130_fd_sc_hd__xor2_1
XFILLER_37_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18333_ _02030_ _02029_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__and2b_1
X_15545_ _08180_ _08189_ vssd1 vssd1 vccd1 vccd1 _08190_ sky130_fd_sc_hd__nor2_1
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _03929_ _05503_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__nor2_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ rbzero.debug_overlay.facingY\[-7\] _04455_ _04482_ _04486_ vssd1 vssd1 vccd1
+ vccd1 _04487_ sky130_fd_sc_hd__a211o_1
XFILLER_72_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18264_ _01951_ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__xnor2_1
X_15476_ _08012_ _08026_ _08119_ vssd1 vssd1 vccd1 vccd1 _08121_ sky130_fd_sc_hd__nand3_1
X_12688_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__and2_1
XFILLER_187_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14427_ _07139_ _07163_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__or2_1
X_17215_ rbzero.wall_tracer.mapX\[9\] _05525_ _09791_ vssd1 vssd1 vccd1 vccd1 _09796_
+ sky130_fd_sc_hd__o21a_1
X_11639_ _04415_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__nor2_1
X_18195_ _01894_ _01895_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__xnor2_1
XFILLER_196_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14358_ _07093_ _07094_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__nor2_2
X_17146_ _07555_ _09763_ rbzero.row_render.size\[8\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00536_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_143_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13309_ _06041_ _06045_ _05991_ _05978_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__or4_1
X_17077_ _09714_ _09716_ vssd1 vssd1 vccd1 vccd1 _09717_ sky130_fd_sc_hd__xor2_4
X_14289_ _07023_ _07025_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__xor2_2
XFILLER_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16028_ _08617_ _08672_ vssd1 vssd1 vccd1 vccd1 _08673_ sky130_fd_sc_hd__nor2_1
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17979_ _01678_ _01679_ _01680_ _09889_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__o31a_1
XFILLER_78_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19718_ _03086_ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20990_ clknet_leaf_14_i_clk _00759_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_38_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03318_ _03318_ vssd1 vssd1 vccd1 vccd1 clknet_0__03318_ sky130_fd_sc_hd__clkbuf_16
X_19649_ _03050_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21611_ net128 _01380_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21542_ net463 _01311_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21473_ net394 _01242_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20424_ rbzero.traced_texa\[-10\] rbzero.texV\[-10\] vssd1 vssd1 vccd1 vccd1 _03334_
+ sky130_fd_sc_hd__nor2_1
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03040_ clknet_0__03040_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03040_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_135_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11990_ _04763_ _04764_ _04345_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__mux2_1
XFILLER_21_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10941_ rbzero.tex_b1\[21\] rbzero.tex_b1\[22\] _03817_ vssd1 vssd1 vccd1 vccd1 _03818_
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13660_ _06363_ _06364_ _06360_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10872_ _03781_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20242__262 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__inv_2
XFILLER_32_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _05346_ _05349_ _05361_ _05364_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__or4_1
XFILLER_25_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _06324_ _06326_ _06327_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__a21oi_1
XFILLER_169_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _07925_ rbzero.wall_tracer.stepDistY\[-2\] vssd1 vssd1 vccd1 vccd1 _07975_
+ sky130_fd_sc_hd__nor2_1
XFILLER_197_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] vssd1
+ vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__xor2_1
XFILLER_197_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15261_ rbzero.debug_overlay.playerY\[-6\] _07905_ vssd1 vssd1 vccd1 vccd1 _07906_
+ sky130_fd_sc_hd__or2_1
XFILLER_185_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12473_ rbzero.wall_tracer.trackDistY\[9\] _05215_ _05217_ rbzero.wall_tracer.trackDistY\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__o22a_1
Xclkbuf_1_0__f__03307_ clknet_0__03307_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03307_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_200_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17000_ _09521_ _09525_ vssd1 vssd1 vccd1 vccd1 _09640_ sky130_fd_sc_hd__nand2_1
XFILLER_126_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14212_ _06947_ _06948_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__or2b_1
X_11424_ _04146_ _04203_ rbzero.row_render.vinf vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15192_ _07841_ _07842_ _07843_ _07844_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__o211ai_2
XFILLER_125_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_8 _07524_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _06857_ _06878_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__nor2_1
XFILLER_67_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11355_ _04088_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__clkbuf_4
XFILLER_193_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _03474_ _03475_ _03478_ _03480_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__and4_1
X_14074_ _06803_ _06810_ vssd1 vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__xor2_1
X_18951_ _02594_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__clkbuf_4
XFILLER_152_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11286_ rbzero.traced_texVinit\[5\] rbzero.spi_registers.vshift\[2\] vssd1 vssd1
+ vccd1 vccd1 _04066_ sky130_fd_sc_hd__or2_1
XFILLER_134_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17902_ _01602_ _01603_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__and2_1
X_13025_ _05605_ _05604_ _05680_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__mux2_1
XFILLER_121_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18882_ _02553_ _02390_ rbzero.wall_tracer.trackDistY\[11\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00624_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_126_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17833_ _10254_ _10276_ _01536_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__a21boi_2
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17764_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__nor2_1
XFILLER_48_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19613__67 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__inv_2
X_14976_ rbzero.wall_tracer.stepDistX\[-5\] _07650_ vssd1 vssd1 vccd1 vccd1 _07658_
+ sky130_fd_sc_hd__nor2_1
X_20325__337 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__inv_2
XFILLER_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19503_ _02980_ _02981_ _02961_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a21o_1
X_16715_ _08062_ _09217_ vssd1 vssd1 vccd1 vccd1 _09357_ sky130_fd_sc_hd__nor2_1
X_13927_ _06031_ _06663_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__nor2_2
X_17695_ _10255_ _10259_ vssd1 vssd1 vccd1 vccd1 _10260_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19434_ _02899_ _02914_ _02915_ _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a31o_1
X_16646_ _08215_ _08985_ _09138_ _08519_ vssd1 vssd1 vccd1 vccd1 _09289_ sky130_fd_sc_hd__o22ai_1
X_13858_ _06564_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__nand2_2
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19365_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__or2_1
X_12809_ rbzero.wall_tracer.mapY\[9\] _05404_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__nor2_1
XFILLER_76_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16577_ _09161_ _09219_ vssd1 vssd1 vccd1 vccd1 _09220_ sky130_fd_sc_hd__nand2_1
XFILLER_188_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13789_ _06520_ _06521_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__nor2_1
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18316_ _09889_ _02015_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__or2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15528_ _07894_ _05490_ vssd1 vssd1 vccd1 vccd1 _08173_ sky130_fd_sc_hd__nand2_1
XFILLER_188_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19296_ rbzero.spi_registers.new_other\[2\] rbzero.spi_registers.spi_buffer\[2\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__mux2_1
XFILLER_188_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18247_ _01943_ _01945_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__nand2_1
XFILLER_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15459_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08104_ sky130_fd_sc_hd__or2_4
XFILLER_176_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18178_ _08895_ _07916_ _07921_ _10134_ _01878_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__o311a_1
XFILLER_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17129_ _09759_ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20070__107 clknet_1_0__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__inv_2
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_1_i_clk clknet_1_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0_1_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_170_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20973_ clknet_leaf_15_i_clk _00742_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21525_ net446 _01294_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21456_ net377 _01225_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21387_ net308 _01156_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__clkinv_2
X_20338_ clknet_1_0__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__buf_1
XFILLER_123_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput56 net56 vssd1 vssd1 vccd1 vccd1 o_gpout[3] sky130_fd_sc_hd__clkbuf_1
XFILLER_150_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput67 net67 vssd1 vssd1 vccd1 vccd1 o_tex_csb sky130_fd_sc_hd__buf_2
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ _03885_ vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14830_ _07486_ _07455_ _07554_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__a21boi_4
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14761_ _07473_ _07477_ _07493_ _07494_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__a31o_1
X_11973_ _04746_ _04747_ _04218_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__mux2_1
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20166__193 clknet_1_1__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__inv_2
XFILLER_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _09140_ _09143_ vssd1 vssd1 vccd1 vccd1 _09144_ sky130_fd_sc_hd__xnor2_2
XFILLER_205_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _06057_ _05982_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__nor2_1
X_10924_ rbzero.tex_b1\[29\] rbzero.tex_b1\[30\] _03806_ vssd1 vssd1 vccd1 vccd1 _03809_
+ sky130_fd_sc_hd__mux2_1
X_17480_ _09952_ _10040_ _10044_ vssd1 vssd1 vccd1 vccd1 _10046_ sky130_fd_sc_hd__and3_1
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14692_ _07379_ _07380_ _05931_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__a21o_1
XFILLER_205_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16431_ _08549_ _08957_ vssd1 vssd1 vccd1 vccd1 _09076_ sky130_fd_sc_hd__xor2_4
X_10855_ _03772_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__clkbuf_1
X_13643_ _06340_ _06342_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19150_ rbzero.otherx\[1\] _02710_ _02715_ _02714_ vssd1 vssd1 vccd1 vccd1 _00730_
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16362_ _08823_ _08059_ _09005_ vssd1 vssd1 vccd1 vccd1 _09007_ sky130_fd_sc_hd__o21ai_1
X_13574_ _05920_ _06016_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__or2_1
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10786_ _03736_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__clkbuf_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _01781_ _01783_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__or2_1
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15313_ _07945_ _07950_ _07956_ _07957_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__a22o_4
X_12525_ _03968_ _03998_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__nor2_1
XFILLER_201_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19081_ rbzero.pov.spi_buffer\[71\] rbzero.pov.ready_buffer\[71\] _02594_ vssd1 vssd1
+ vccd1 vccd1 _02673_ sky130_fd_sc_hd__mux2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16293_ _08806_ _08801_ _08805_ vssd1 vssd1 vccd1 vccd1 _08938_ sky130_fd_sc_hd__a21bo_1
XFILLER_121_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18032_ _01626_ _01628_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__nor2_1
XFILLER_200_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12456_ _05210_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__buf_6
XFILLER_157_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15244_ rbzero.wall_tracer.wall\[1\] _03999_ _05280_ _03996_ vssd1 vssd1 vccd1 vccd1
+ _07891_ sky130_fd_sc_hd__a22o_1
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11407_ rbzero.row_render.size\[4\] _04150_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__xnor2_1
X_15175_ _07816_ _07824_ _07828_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__a21oi_1
X_12387_ _03474_ _04814_ _04317_ _04809_ _05146_ _05145_ vssd1 vssd1 vccd1 vccd1 _05154_
+ sky130_fd_sc_hd__mux4_1
XFILLER_158_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14126_ _06827_ _06829_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ _04097_ _04114_ _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__or3_1
X_19983_ rbzero.pov.ready_buffer\[32\] _03247_ _03249_ rbzero.debug_overlay.facingY\[10\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__a221o_1
XFILLER_180_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14057_ _06789_ _06793_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__xnor2_1
X_18934_ _02596_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11269_ rbzero.traced_texVinit\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _04049_
+ sky130_fd_sc_hd__nand2_1
XFILLER_141_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13008_ _05642_ _05744_ _05634_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a21oi_1
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18865_ _02530_ _02532_ _02531_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__o21bai_1
XFILLER_122_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17816_ _09114_ _09693_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__nor2_1
XFILLER_39_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18796_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.stepDistY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__nand2_1
XFILLER_43_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17747_ _01443_ _01444_ _01450_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__a21oi_1
XFILLER_94_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14959_ rbzero.wall_tracer.trackDistX\[11\] rbzero.wall_tracer.trackDistY\[11\] _04019_
+ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__a21o_1
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17678_ _10241_ _10242_ vssd1 vssd1 vccd1 vccd1 _10243_ sky130_fd_sc_hd__xnor2_2
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19417_ _02885_ _02901_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16629_ _09114_ _08204_ vssd1 vssd1 vccd1 vccd1 _09272_ sky130_fd_sc_hd__nor2_1
XFILLER_126_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19348_ rbzero.debug_overlay.vplaneY\[-9\] _07703_ _07855_ rbzero.wall_tracer.rayAddendY\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a22o_1
XFILLER_149_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19279_ _02794_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21310_ net231 _01079_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_176_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21241_ clknet_leaf_87_i_clk _01010_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21172_ clknet_leaf_78_i_clk _00941_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20054_ rbzero.spi_registers.got_new_vinf _09753_ _02728_ _02555_ vssd1 vssd1 vccd1
+ vccd1 _01061_ sky130_fd_sc_hd__a31o_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20308__321 clknet_1_0__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__inv_2
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20956_ clknet_leaf_99_i_clk _00725_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20887_ clknet_leaf_87_i_clk _00656_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10640_ rbzero.tex_g1\[36\] rbzero.tex_g1\[37\] _03658_ vssd1 vssd1 vccd1 vccd1 _03660_
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _03613_ vssd1 vssd1 vccd1 vccd1 _03623_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12310_ _05034_ net25 _05051_ _05061_ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__a311o_2
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21508_ net429 _01277_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13290_ _05855_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__xnor2_1
XFILLER_177_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20354__363 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__inv_2
XFILLER_5_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12241_ net19 _04996_ _05010_ _04867_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__or4b_1
XFILLER_181_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21439_ net360 _01208_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12172_ _04813_ _04811_ _04006_ _03475_ _04910_ net9 vssd1 vssd1 vccd1 vccd1 _04943_
+ sky130_fd_sc_hd__mux4_1
XFILLER_135_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11123_ net71 _03480_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__nand2_4
XFILLER_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16980_ _08160_ _09483_ vssd1 vssd1 vccd1 vccd1 _09620_ sky130_fd_sc_hd__nor2_1
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15931_ _08573_ _08575_ vssd1 vssd1 vccd1 vccd1 _08576_ sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_64_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11054_ rbzero.tex_b0\[32\] rbzero.tex_b0\[31\] _03876_ vssd1 vssd1 vccd1 vccd1 _03877_
+ sky130_fd_sc_hd__mux2_1
XFILLER_153_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18650_ _01739_ _09162_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__nor2_1
XFILLER_190_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _08152_ _08153_ vssd1 vssd1 vccd1 vccd1 _08507_ sky130_fd_sc_hd__nand2_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17601_ _10165_ _10166_ vssd1 vssd1 vccd1 vccd1 _10167_ sky130_fd_sc_hd__or2b_1
XFILLER_18_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14813_ rbzero.wall_tracer.stepDistY\[-4\] _07541_ _07461_ vssd1 vssd1 vccd1 vccd1
+ _07542_ sky130_fd_sc_hd__mux2_1
XFILLER_92_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ _02272_ _02277_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__and2_1
XFILLER_149_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _08413_ _08437_ vssd1 vssd1 vccd1 vccd1 _08438_ sky130_fd_sc_hd__xnor2_2
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_102 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_102/HI zeros[12]
+ sky130_fd_sc_hd__conb_1
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17532_ _10096_ _10097_ vssd1 vssd1 vccd1 vccd1 _10098_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_79_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_i_clk
+ sky130_fd_sc_hd__clkbuf_16
Xtop_ew_algofoogle_113 vssd1 vssd1 vccd1 vccd1 ones[7] top_ew_algofoogle_113/LO sky130_fd_sc_hd__conb_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14744_ _07385_ _07387_ vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__or2b_1
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _04726_ _04728_ _04731_ _04332_ _04241_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__a221o_1
XFILLER_189_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ rbzero.tex_b1\[37\] rbzero.tex_b1\[38\] _03795_ vssd1 vssd1 vccd1 vccd1 _03800_
+ sky130_fd_sc_hd__mux2_1
X_17463_ rbzero.wall_tracer.trackDistX\[0\] rbzero.wall_tracer.stepDistX\[0\] vssd1
+ vssd1 vccd1 vccd1 _10030_ sky130_fd_sc_hd__nor2_1
X_14675_ _06724_ _06761_ _07411_ _07340_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__o211a_1
X_11887_ rbzero.color_sky\[3\] rbzero.color_floor\[3\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04664_ sky130_fd_sc_hd__mux2_1
X_19202_ rbzero.spi_registers.new_sky\[4\] rbzero.spi_registers.got_new_sky _02711_
+ _02741_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__a31o_1
XFILLER_189_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16414_ _09056_ _09058_ vssd1 vssd1 vccd1 vccd1 _09059_ sky130_fd_sc_hd__xnor2_2
XFILLER_177_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13626_ _06361_ _06362_ _06078_ _05982_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a211o_1
X_10838_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _03762_ vssd1 vssd1 vccd1 vccd1 _03764_
+ sky130_fd_sc_hd__mux2_1
X_17394_ _09661_ _08356_ _09960_ vssd1 vssd1 vccd1 vccd1 _09961_ sky130_fd_sc_hd__or3_1
XFILLER_125_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19133_ _02701_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16345_ _08987_ _08989_ vssd1 vssd1 vccd1 vccd1 _08990_ sky130_fd_sc_hd__xnor2_2
X_10769_ _03727_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__clkbuf_1
X_13557_ _05995_ _06113_ _06045_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__a21o_1
XFILLER_160_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19064_ _02664_ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__clkbuf_1
X_12508_ rbzero.wall_tracer.trackDistX\[-4\] vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__inv_2
X_16276_ _08869_ _08919_ vssd1 vssd1 vccd1 vccd1 _08921_ sky130_fd_sc_hd__or2_1
XFILLER_121_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13488_ _06197_ _06198_ _06224_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__o21ai_1
XFILLER_201_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18015_ _01616_ _01617_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__nand2_1
X_15227_ rbzero.wall_tracer.rayAddendX\[9\] _00013_ _07831_ _07875_ _07877_ vssd1
+ vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_17_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12439_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__buf_6
XFILLER_201_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15158_ _07800_ _07812_ vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__xor2_1
XFILLER_141_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14109_ _06763_ _06845_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__xnor2_2
XFILLER_141_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15089_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.debug_overlay.vplaneX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _07749_ sky130_fd_sc_hd__nor2_1
X_19966_ rbzero.pov.ready_buffer\[39\] _03247_ _03249_ rbzero.debug_overlay.facingX\[-3\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__a221o_1
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18917_ rbzero.spi_registers.spi_counter\[3\] _02580_ vssd1 vssd1 vccd1 vccd1 _02584_
+ sky130_fd_sc_hd__or2_1
XFILLER_132_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19897_ rbzero.pov.ready_buffer\[46\] _02823_ _03193_ _03201_ vssd1 vssd1 vccd1 vccd1
+ _03202_ sky130_fd_sc_hd__a211o_1
XFILLER_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18848_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.stepDistY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__or2_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20182__208 clknet_1_0__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__inv_2
X_18779_ _09812_ _09597_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__nand2_1
X_20810_ clknet_leaf_66_i_clk _00579_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20741_ clknet_leaf_71_i_clk _00510_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.side
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20672_ clknet_leaf_60_i_clk _00456_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_149_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21224_ clknet_leaf_24_i_clk _00993_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21155_ clknet_leaf_68_i_clk _00924_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21086_ net176 _00855_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20037_ _03277_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__clkbuf_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _04582_ _04584_ _04587_ _04208_ _04142_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__a221o_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _05532_ _05283_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__nor2_4
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _03478_ _04026_ _04047_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a21oi_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20939_ clknet_leaf_9_i_clk _00708_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _07170_ _07182_ _07196_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__o21ai_1
X_11672_ _04004_ _04419_ _04450_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__and3b_1
XFILLER_183_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10623_ rbzero.tex_g1\[44\] rbzero.tex_g1\[45\] _03647_ vssd1 vssd1 vccd1 vccd1 _03651_
+ sky130_fd_sc_hd__mux2_1
X_13411_ _06144_ _06091_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__xnor2_1
X_14391_ _06675_ _06761_ _07108_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__o21ai_1
XFILLER_168_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20278__294 clknet_1_0__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__inv_2
XFILLER_31_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16130_ _08773_ _08772_ vssd1 vssd1 vccd1 vccd1 _08775_ sky130_fd_sc_hd__or2b_1
XFILLER_127_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13342_ _06053_ _06056_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__and2_1
X_10554_ _03614_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13273_ _05973_ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__nor2_1
X_16061_ _08594_ _08705_ vssd1 vssd1 vccd1 vccd1 _08706_ sky130_fd_sc_hd__nor2_1
X_10485_ rbzero.tex_r0\[46\] rbzero.tex_r0\[45\] _03569_ vssd1 vssd1 vccd1 vccd1 _03578_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12224_ _04987_ _04988_ _04991_ _04993_ net16 _04960_ vssd1 vssd1 vccd1 vccd1 _04994_
+ sky130_fd_sc_hd__mux4_1
XFILLER_170_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15012_ rbzero.wall_tracer.state\[14\] _04037_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__nand2_2
XFILLER_135_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19820_ _03140_ rbzero.pov.ready_buffer\[59\] _03141_ vssd1 vssd1 vccd1 vccd1 _03142_
+ sky130_fd_sc_hd__mux2_1
X_12155_ net51 _04904_ net47 vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__a21o_1
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11106_ rbzero.tex_b0\[7\] rbzero.tex_b0\[6\] _03898_ vssd1 vssd1 vccd1 vccd1 _03904_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__03320_ clknet_0__03320_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03320_
+ sky130_fd_sc_hd__clkbuf_16
X_19751_ rbzero.pov.spi_buffer\[49\] rbzero.pov.spi_buffer\[50\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03104_ sky130_fd_sc_hd__mux2_1
XFILLER_110_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12086_ net43 _04857_ _04838_ net41 vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__a22o_1
XFILLER_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16963_ _09085_ _09603_ vssd1 vssd1 vccd1 vccd1 _09604_ sky130_fd_sc_hd__nand2_1
XFILLER_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18702_ _09808_ _02396_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__nand2_1
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15914_ _07923_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08559_ sky130_fd_sc_hd__or3_1
XFILLER_77_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11037_ rbzero.tex_b0\[40\] rbzero.tex_b0\[39\] _03865_ vssd1 vssd1 vccd1 vccd1 _03868_
+ sky130_fd_sc_hd__mux2_1
X_19682_ _03067_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__clkbuf_1
X_16894_ _09533_ _09534_ vssd1 vssd1 vccd1 vccd1 _09535_ sky130_fd_sc_hd__xor2_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18633_ _02327_ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__xnor2_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15845_ _07945_ rbzero.wall_tracer.stepDistX\[-11\] vssd1 vssd1 vccd1 vccd1 _08490_
+ sky130_fd_sc_hd__nand2_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18564_ _01739_ _09027_ _02260_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__or3_1
XFILLER_40_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15776_ _08062_ _08158_ _08150_ _08054_ vssd1 vssd1 vccd1 vccd1 _08421_ sky130_fd_sc_hd__o22a_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12988_ _05665_ _05666_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__nand2_1
XFILLER_75_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17515_ _09664_ _09665_ _09945_ vssd1 vssd1 vccd1 vccd1 _10081_ sky130_fd_sc_hd__a21oi_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14727_ _05892_ _07395_ _07398_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__o21a_1
X_19583__39 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__inv_2
XFILLER_205_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18495_ _02185_ _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__xor2_1
X_11939_ _04712_ _04713_ _04714_ _04247_ _04306_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__o221a_1
XFILLER_75_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17446_ _09680_ _09721_ _10012_ vssd1 vssd1 vccd1 vccd1 _10013_ sky130_fd_sc_hd__a21o_1
X_14658_ _07352_ _07362_ _05779_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ _06281_ _06283_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17377_ _09245_ _08427_ vssd1 vssd1 vccd1 vccd1 _09944_ sky130_fd_sc_hd__nor2_1
XFILLER_158_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14589_ _07131_ _07325_ _07206_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__a21oi_1
XFILLER_174_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19116_ _02692_ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16328_ _07981_ _07989_ _08189_ _08971_ vssd1 vssd1 vccd1 vccd1 _08973_ sky130_fd_sc_hd__or4_1
XFILLER_185_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19047_ _02655_ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16259_ _08892_ _08899_ _08903_ vssd1 vssd1 vccd1 vccd1 _08904_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19949_ rbzero.pov.ready _02707_ _02820_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__and3_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20724_ clknet_leaf_82_i_clk _00493_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_24_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_6_0_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20655_ clknet_leaf_52_i_clk _00439_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20586_ rbzero.wall_tracer.rayAddendX\[-7\] _03443_ _07756_ _03455_ vssd1 vssd1 vccd1
+ vccd1 _01426_ sky130_fd_sc_hd__a22o_1
XFILLER_164_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21207_ clknet_leaf_28_i_clk _00976_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21138_ clknet_leaf_97_i_clk _00907_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13960_ _06696_ _06671_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__nor2_1
XFILLER_47_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21069_ net159 _00838_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12911_ _05646_ _05647_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__xnor2_4
XFILLER_207_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13891_ _06572_ _06627_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ _07951_ rbzero.wall_tracer.stepDistY\[-1\] _08272_ _08274_ vssd1 vssd1 vccd1
+ vccd1 _08275_ sky130_fd_sc_hd__a22oi_4
X_12842_ _04030_ _05346_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__a21o_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _08193_ _08205_ vssd1 vssd1 vccd1 vccd1 _08206_ sky130_fd_sc_hd__xnor2_4
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _05518_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__clkbuf_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _09871_ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _07247_ _07248_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__nor2_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _01882_ _01877_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__and2b_1
XFILLER_159_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ rbzero.debug_overlay.playerY\[0\] _04459_ _04460_ rbzero.debug_overlay.playerY\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__a22o_1
X_15492_ _08131_ _08136_ vssd1 vssd1 vccd1 vccd1 _08137_ sky130_fd_sc_hd__xor2_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.stepDistX\[-12\]
+ _09809_ vssd1 vssd1 vccd1 vccd1 _09810_ sky130_fd_sc_hd__a21o_1
X_14443_ _07176_ _07178_ _07179_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11655_ gpout0.hpos\[6\] _04430_ _04431_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__and3_1
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10606_ _03641_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17162_ _07706_ vssd1 vssd1 vccd1 vccd1 _09768_ sky130_fd_sc_hd__clkbuf_4
X_11586_ rbzero.tex_r1\[25\] rbzero.tex_r1\[24\] _04342_ vssd1 vssd1 vccd1 vccd1 _04365_
+ sky130_fd_sc_hd__mux2_1
X_14374_ _06689_ _07072_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__nor2_1
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16113_ _08737_ _08757_ vssd1 vssd1 vccd1 vccd1 _08758_ sky130_fd_sc_hd__nor2_1
X_10537_ _03605_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13325_ _06059_ _06060_ _06061_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__a21oi_2
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17093_ _09730_ _09732_ vssd1 vssd1 vccd1 vccd1 _09733_ sky130_fd_sc_hd__xor2_2
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16044_ _08683_ _08688_ vssd1 vssd1 vccd1 vccd1 _08689_ sky130_fd_sc_hd__or2b_1
X_10468_ _03557_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__clkbuf_4
X_13256_ _05988_ _05989_ _05992_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__and3_1
XFILLER_170_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12207_ net17 vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__inv_2
XFILLER_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13187_ _05695_ _05724_ _05793_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__mux2_1
X_10399_ rbzero.tex_r1\[20\] rbzero.tex_r1\[21\] _03527_ vssd1 vssd1 vccd1 vccd1 _03531_
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12138_ net8 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__inv_2
X_19803_ _03130_ vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__clkbuf_1
X_17995_ _01566_ _01696_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__xnor2_1
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03303_ clknet_0__03303_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03303_
+ sky130_fd_sc_hd__clkbuf_16
X_12069_ _04840_ net61 vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__or2_1
X_16946_ _09476_ _09586_ vssd1 vssd1 vccd1 vccd1 _09587_ sky130_fd_sc_hd__xnor2_1
X_19734_ rbzero.pov.spi_buffer\[41\] rbzero.pov.spi_buffer\[42\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03095_ sky130_fd_sc_hd__mux2_1
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19665_ _03058_ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16877_ _09393_ _09402_ _09400_ vssd1 vssd1 vccd1 vccd1 _09518_ sky130_fd_sc_hd__a21o_1
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18616_ _02125_ _02128_ _02222_ _02223_ _02312_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__a311oi_2
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _07995_ _07981_ _07989_ _07931_ vssd1 vssd1 vccd1 vccd1 _08473_ sky130_fd_sc_hd__o22ai_2
XFILLER_93_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18547_ _02151_ _02243_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__xnor2_1
X_15759_ _08396_ _08392_ vssd1 vssd1 vccd1 vccd1 _08404_ sky130_fd_sc_hd__or2b_1
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18478_ _02174_ _02175_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__nand2_1
XFILLER_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17429_ _08519_ _09699_ vssd1 vssd1 vccd1 vccd1 _09996_ sky130_fd_sc_hd__or2_1
XFILLER_53_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20440_ _03272_ _03346_ _03347_ _03327_ rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1
+ _01388_ sky130_fd_sc_hd__a32o_1
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20371_ clknet_1_0__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__buf_1
XFILLER_173_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20707_ clknet_leaf_73_i_clk _00013_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11440_ _04215_ _04216_ _04219_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
XFILLER_138_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20638_ clknet_leaf_65_i_clk _00422_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11371_ rbzero.row_render.size\[5\] rbzero.row_render.size\[4\] _04150_ vssd1 vssd1
+ vccd1 vccd1 _04151_ sky130_fd_sc_hd__or3_1
X_20569_ gpout0.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__nor2_1
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ _03490_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13110_ _05798_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__inv_2
X_14090_ _06805_ _06740_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__nor2_1
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13041_ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__clkbuf_4
XFILLER_180_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16800_ _09415_ _09441_ vssd1 vssd1 vccd1 vccd1 _09442_ sky130_fd_sc_hd__xnor2_2
X_17780_ _01482_ _01483_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__and2b_1
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14992_ _07666_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16731_ _09092_ _09095_ _09229_ vssd1 vssd1 vccd1 vccd1 _09373_ sky130_fd_sc_hd__a21oi_1
XFILLER_87_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13943_ _06161_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__clkbuf_4
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19450_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.debug_overlay.vplaneY\[-6\] _02930_
+ _02931_ _03913_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__o41a_1
X_16662_ _09275_ _09303_ _09304_ vssd1 vssd1 vccd1 vccd1 _09305_ sky130_fd_sc_hd__nand3_1
X_13874_ _06607_ _06610_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__and2b_1
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18401_ _02065_ _02099_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__xor2_1
X_15613_ _08257_ _08238_ vssd1 vssd1 vccd1 vccd1 _08258_ sky130_fd_sc_hd__nor2_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12825_ _05561_ _05492_ _05493_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__or3_2
X_19381_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__or2_1
XFILLER_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16593_ _09234_ _09235_ vssd1 vssd1 vccd1 vccd1 _09236_ sky130_fd_sc_hd__nor2_1
XFILLER_90_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18332_ _02029_ _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__and2b_1
XFILLER_91_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15544_ _08147_ rbzero.wall_tracer.stepDistX\[2\] _08188_ vssd1 vssd1 vccd1 vccd1
+ _08189_ sky130_fd_sc_hd__a21boi_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12756_ _05496_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__inv_2
XFILLER_203_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18263_ _01960_ _01962_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__xor2_1
XFILLER_124_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ rbzero.debug_overlay.facingY\[-8\] _04466_ _04483_ _04485_ vssd1 vssd1 vccd1
+ vccd1 _04486_ sky130_fd_sc_hd__a211o_1
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15475_ _08012_ _08026_ _08119_ vssd1 vssd1 vccd1 vccd1 _08120_ sky130_fd_sc_hd__a21o_1
X_12687_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] _05434_
+ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__and3_1
XFILLER_147_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17214_ rbzero.wall_tracer.mapX\[9\] _09781_ _09779_ _09795_ vssd1 vssd1 vccd1 vccd1
+ _00574_ sky130_fd_sc_hd__a22o_1
X_14426_ _06724_ _06663_ _07138_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__o21a_1
X_18194_ _01770_ _01771_ _01772_ _01775_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a31o_1
X_11638_ _04024_ _04416_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__or2_2
XFILLER_200_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17145_ _07552_ _09763_ rbzero.row_render.size\[7\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00535_ sky130_fd_sc_hd__a2bb2o_1
X_14357_ _07090_ _07092_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__and2_1
XFILLER_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11569_ _04136_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__buf_4
XFILLER_156_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13308_ _05899_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__clkbuf_4
X_20137__168 clknet_1_0__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__inv_2
XFILLER_170_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17076_ _09559_ _09570_ _09715_ vssd1 vssd1 vccd1 vccd1 _09716_ sky130_fd_sc_hd__a21oi_2
XFILLER_115_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14288_ _06757_ _06797_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__a21boi_2
XFILLER_157_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16027_ _08619_ _08671_ vssd1 vssd1 vccd1 vccd1 _08672_ sky130_fd_sc_hd__and2b_1
X_13239_ _05974_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__nor2_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17978_ _01678_ _01679_ _01680_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__o21ai_1
X_16929_ _09567_ _09569_ vssd1 vssd1 vccd1 vccd1 _09570_ sky130_fd_sc_hd__xor2_2
X_19717_ rbzero.pov.spi_buffer\[33\] rbzero.pov.spi_buffer\[34\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03086_ sky130_fd_sc_hd__mux2_1
XFILLER_168_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03317_ _03317_ vssd1 vssd1 vccd1 vccd1 clknet_0__03317_ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19648_ rbzero.pov.spi_buffer\[0\] rbzero.pov.spi_buffer\[1\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03050_ sky130_fd_sc_hd__mux2_1
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20302__316 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__inv_2
X_21610_ net127 _01379_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21541_ net462 _01310_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21472_ net393 _01241_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20423_ _03329_ _03330_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__and2_1
XFILLER_135_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_11_0_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_11_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10940_ _03646_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__clkbuf_4
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ rbzero.tex_b1\[54\] rbzero.tex_b1\[55\] _03773_ vssd1 vssd1 vccd1 vccd1 _03781_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _05362_ _05363_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__and2_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13590_ _06304_ _06323_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__nor2_1
XFILLER_197_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12541_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] _05290_
+ _05293_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__a221o_2
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_i_clk clknet_1_1_1_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__or3_1
XFILLER_71_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__03306_ clknet_0__03306_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03306_
+ sky130_fd_sc_hd__clkbuf_16
X_12472_ _05221_ _05226_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__nor2_1
X_14211_ _06932_ _06945_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__xnor2_1
XFILLER_71_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11423_ rbzero.row_render.size\[10\] rbzero.row_render.size\[9\] _04153_ _04202_
+ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__or4_1
XFILLER_172_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15191_ _07785_ rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 _07844_
+ sky130_fd_sc_hd__or2_1
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 _07530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14142_ _06857_ _06878_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__xor2_1
X_11354_ rbzero.floor_leak\[4\] _04121_ _04116_ rbzero.floor_leak\[5\] vssd1 vssd1
+ vccd1 vccd1 _04134_ sky130_fd_sc_hd__o22a_1
XFILLER_67_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10305_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__buf_6
XFILLER_180_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18950_ _02604_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__clkbuf_1
X_14073_ _06776_ _06740_ _06804_ _06809_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__o31a_1
XFILLER_4_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11285_ rbzero.texV\[6\] _04064_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__xor2_1
XFILLER_140_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17901_ _01602_ _01603_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__nor2_1
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13024_ _05677_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__inv_2
XFILLER_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18881_ _05532_ _02552_ _02399_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__o21a_1
X_17832_ _10273_ _10275_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__or2b_1
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17763_ _09249_ _09359_ _10206_ _10205_ _09391_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__o32a_1
XFILLER_48_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14975_ _00008_ _07530_ _07657_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16714_ _09354_ _09355_ vssd1 vssd1 vccd1 vccd1 _09356_ sky130_fd_sc_hd__xnor2_1
X_19502_ _02905_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 _02981_
+ sky130_fd_sc_hd__nand2_1
XFILLER_207_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13926_ _06662_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__clkbuf_4
X_17694_ _09292_ _09695_ _08895_ vssd1 vssd1 vccd1 vccd1 _10259_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19433_ _03912_ _02916_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__nand2_1
XFILLER_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16645_ _09284_ _09287_ _05210_ vssd1 vssd1 vccd1 vccd1 _09288_ sky130_fd_sc_hd__a21o_1
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857_ _06273_ _06593_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__xor2_1
XFILLER_179_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19364_ _02851_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__or2b_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12808_ rbzero.wall_tracer.mapY\[9\] _05404_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__and2_1
X_16576_ _09214_ _09218_ vssd1 vssd1 vccd1 vccd1 _09219_ sky130_fd_sc_hd__xnor2_1
X_13788_ _06507_ _06523_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__nand2_1
X_18315_ _02013_ _02014_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__xnor2_1
XFILLER_163_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ _07560_ _08171_ vssd1 vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__xnor2_1
X_12739_ _05440_ _05465_ _05462_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__a21boi_1
X_19295_ _02803_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__clkbuf_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18246_ _01943_ _01945_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__or2_1
XFILLER_148_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15458_ _05197_ rbzero.wall_tracer.stepDistX\[-8\] vssd1 vssd1 vccd1 vccd1 _08103_
+ sky130_fd_sc_hd__nor2_2
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14409_ _06239_ _07111_ _07145_ _07131_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__o31a_1
X_18177_ _08895_ _08767_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__nand2_1
XFILLER_204_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ _07990_ _05496_ _08028_ _08033_ vssd1 vssd1 vccd1 vccd1 _08034_ sky130_fd_sc_hd__o31a_4
XFILLER_190_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17128_ _04446_ _09750_ _09758_ vssd1 vssd1 vccd1 vccd1 _09759_ sky130_fd_sc_hd__and3_1
XFILLER_144_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17059_ _09283_ rbzero.wall_tracer.stepDistY\[11\] _08235_ _09698_ vssd1 vssd1 vccd1
+ vccd1 _09699_ sky130_fd_sc_hd__a22oi_4
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20972_ clknet_leaf_15_i_clk _00741_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21524_ net445 _01293_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21455_ net376 _01224_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21386_ net307 _01155_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput57 net57 vssd1 vssd1 vccd1 vccd1 o_gpout[4] sky130_fd_sc_hd__clkbuf_1
XFILLER_134_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11070_ rbzero.tex_b0\[24\] rbzero.tex_b0\[23\] _03876_ vssd1 vssd1 vccd1 vccd1 _03885_
+ sky130_fd_sc_hd__mux2_1
Xoutput68 net68 vssd1 vssd1 vccd1 vccd1 o_tex_oeb0 sky130_fd_sc_hd__buf_2
XFILLER_115_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20056__94 clknet_1_1__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__inv_2
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14760_ _07102_ _05952_ _05844_ _07366_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__and4b_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11972_ rbzero.tex_b1\[25\] rbzero.tex_b1\[24\] _04342_ vssd1 vssd1 vccd1 vccd1 _04747_
+ sky130_fd_sc_hd__mux2_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _06442_ _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__xor2_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _03808_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__clkbuf_1
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _07378_ _07413_ _07414_ _07427_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__o31a_1
XFILLER_186_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16430_ rbzero.debug_overlay.playerY\[-7\] rbzero.debug_overlay.playerX\[-7\] _07895_
+ vssd1 vssd1 vccd1 vccd1 _09075_ sky130_fd_sc_hd__mux2_1
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ _06347_ _06373_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__xnor2_2
X_10854_ rbzero.tex_b1\[62\] rbzero.tex_b1\[63\] _03691_ vssd1 vssd1 vccd1 vccd1 _03772_
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16361_ _08823_ _08058_ _09005_ vssd1 vssd1 vccd1 vccd1 _09006_ sky130_fd_sc_hd__or3_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13573_ _05823_ _05939_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__or2_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ rbzero.tex_g0\[32\] rbzero.tex_g0\[31\] _03729_ vssd1 vssd1 vccd1 vccd1 _03736_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18100_ _01667_ _01800_ _01787_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__a21o_1
XFILLER_158_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15312_ rbzero.wall_tracer.visualWallDist\[-4\] _07925_ _05207_ vssd1 vssd1 vccd1
+ vccd1 _07957_ sky130_fd_sc_hd__a21oi_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19080_ _02672_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__clkbuf_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _05278_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__inv_2
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _08764_ _08807_ vssd1 vssd1 vccd1 vccd1 _08937_ sky130_fd_sc_hd__xor2_1
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18031_ _01698_ _01732_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__xor2_1
XFILLER_201_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15243_ _07890_ vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__clkbuf_1
X_12455_ _05209_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__buf_4
XFILLER_184_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11406_ _04151_ _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__nand2_1
XFILLER_126_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15174_ _07785_ rbzero.wall_tracer.rayAddendX\[6\] vssd1 vssd1 vccd1 vccd1 _07828_
+ sky130_fd_sc_hd__xnor2_1
X_12386_ net35 vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__inv_2
XFILLER_165_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20331__342 clknet_1_0__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__inv_2
X_14125_ _06846_ _06847_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__xor2_2
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11337_ _04096_ _04075_ _04093_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__nor3_1
XFILLER_207_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19982_ net70 _03247_ _03249_ rbzero.debug_overlay.facingY\[0\] _03251_ vssd1 vssd1
+ vccd1 vccd1 _01024_ sky130_fd_sc_hd__a221o_1
XFILLER_98_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14056_ _06787_ _06791_ _06792_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__o21ai_1
X_18933_ rbzero.pov.spi_buffer\[0\] rbzero.pov.ready_buffer\[0\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02596_ sky130_fd_sc_hd__mux2_1
XFILLER_98_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _04048_
+ sky130_fd_sc_hd__nand2_1
XFILLER_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13007_ _05622_ _05635_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__xnor2_2
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18864_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.stepDistY\[9\] vssd1
+ vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__nand2_1
X_11199_ rbzero.map_rom.f4 _03933_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__xnor2_1
X_17815_ _01514_ _01518_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18795_ _02478_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17746_ _01448_ _01449_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__nand2_1
X_14958_ _04019_ _07647_ _07648_ _07642_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__o211a_1
XFILLER_36_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13909_ _05752_ _06201_ _06621_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17677_ _10094_ _08057_ vssd1 vssd1 vccd1 vccd1 _10242_ sky130_fd_sc_hd__nor2_1
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14889_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.trackDistX\[-10\]
+ _07592_ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__mux2_1
XFILLER_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16628_ _09119_ _09270_ vssd1 vssd1 vccd1 vccd1 _09271_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19416_ _02899_ _02900_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__nand2_1
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16559_ rbzero.wall_tracer.texu\[1\] _09085_ vssd1 vssd1 vccd1 vccd1 _09203_ sky130_fd_sc_hd__or2_1
X_19347_ _02826_ _02837_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19278_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_leak\[1\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__mux2_1
XFILLER_176_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18229_ _01838_ _01852_ _01850_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__a21o_1
XFILLER_50_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21240_ clknet_leaf_87_i_clk _01009_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_163_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21171_ clknet_leaf_78_i_clk _00940_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20053_ _03285_ _03288_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__nor2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19589__45 clknet_1_0__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__inv_2
XFILLER_46_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ clknet_leaf_99_i_clk _00724_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ clknet_leaf_87_i_clk _00655_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10570_ _03622_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21507_ net428 _01276_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12240_ _04960_ _04961_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__nand2_1
X_21438_ net359 _01207_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12171_ net11 _04908_ _04937_ _04941_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__a31o_1
X_21369_ net290 _01138_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11122_ _03911_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_8
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15930_ _08498_ _08574_ vssd1 vssd1 vccd1 vccd1 _08575_ sky130_fd_sc_hd__xnor2_1
X_11053_ _03717_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _08489_ _08505_ vssd1 vssd1 vccd1 vccd1 _08506_ sky130_fd_sc_hd__or2b_1
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ _10037_ _10038_ _10164_ vssd1 vssd1 vccd1 vccd1 _10166_ sky130_fd_sc_hd__a21o_1
Xclkbuf_0_i_clk i_clk vssd1 vssd1 vccd1 vccd1 clknet_0_i_clk sky130_fd_sc_hd__clkbuf_16
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ _07486_ _07455_ _07539_ _07527_ _07540_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__a221o_4
XFILLER_92_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18580_ _02275_ _02276_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__xor2_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _08435_ _08436_ vssd1 vssd1 vccd1 vccd1 _08437_ sky130_fd_sc_hd__and2_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ _08275_ _08356_ vssd1 vssd1 vccd1 vccd1 _10097_ sky130_fd_sc_hd__nor2_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_103 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_103/HI zeros[13]
+ sky130_fd_sc_hd__conb_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _07475_ _07476_ _07477_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_114 vssd1 vssd1 vccd1 vccd1 ones[8] top_ew_algofoogle_114/LO sky130_fd_sc_hd__conb_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11955_ _04729_ _04730_ _04329_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__mux2_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ _03799_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__clkbuf_1
X_17462_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _10029_ sky130_fd_sc_hd__nand2_1
X_14674_ _06239_ _07149_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__nor2_1
X_11886_ _04628_ _04206_ _04662_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__or3b_1
X_16413_ _08169_ _08469_ _09057_ vssd1 vssd1 vccd1 vccd1 _09058_ sky130_fd_sc_hd__a21o_1
X_19201_ _02747_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__clkbuf_1
X_13625_ _06041_ _06031_ _06285_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__o21ai_1
X_17393_ _09663_ _09959_ vssd1 vssd1 vccd1 vccd1 _09960_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10837_ _03763_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__clkbuf_1
X_19132_ rbzero.spi_registers.sclk_buffer\[1\] rbzero.spi_registers.sclk_buffer\[0\]
+ _05189_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__mux2_1
X_16344_ _08237_ _08239_ _08229_ _08988_ vssd1 vssd1 vccd1 vccd1 _08989_ sky130_fd_sc_hd__o31a_1
XFILLER_125_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13556_ _06057_ _05940_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__nor2_1
X_10768_ rbzero.tex_g0\[40\] rbzero.tex_g0\[39\] _03718_ vssd1 vssd1 vccd1 vccd1 _03727_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19063_ rbzero.pov.spi_buffer\[62\] rbzero.pov.ready_buffer\[62\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02664_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_12507_ _05258_ rbzero.wall_tracer.trackDistX\[-1\] _05251_ rbzero.wall_tracer.trackDistX\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__a22o_1
X_16275_ _08869_ _08919_ vssd1 vssd1 vccd1 vccd1 _08920_ sky130_fd_sc_hd__nand2_1
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13487_ _06209_ _06223_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__xnor2_1
X_10699_ _03690_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__clkbuf_1
X_18014_ _01474_ _08423_ _01596_ _01594_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__o31a_1
XFILLER_201_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15226_ _07858_ _07862_ _07876_ _04034_ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__a211o_1
XFILLER_173_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12438_ _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__buf_4
XFILLER_201_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15157_ _07785_ _04462_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__xor2_1
X_12369_ _05115_ _05123_ _05130_ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__or4_2
XFILLER_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14108_ _06704_ _06668_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__nor2_1
XFILLER_99_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15088_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.debug_overlay.vplaneX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__and2_1
X_19965_ _02695_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18916_ rbzero.spi_registers.spi_counter\[3\] _02580_ vssd1 vssd1 vccd1 vccd1 _02583_
+ sky130_fd_sc_hd__and2_1
X_14039_ _05984_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__buf_2
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19896_ _08004_ _03141_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__nor2_1
XFILLER_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18847_ _02523_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18778_ _02463_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__clkbuf_1
X_17729_ _10292_ _10293_ vssd1 vssd1 vccd1 vccd1 _10294_ sky130_fd_sc_hd__nor2_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20740_ clknet_leaf_45_i_clk _00509_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.wall\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20671_ clknet_leaf_61_i_clk _00455_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21223_ clknet_leaf_22_i_clk _00992_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_191_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21154_ clknet_leaf_86_i_clk _00923_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20105_ clknet_1_1__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__buf_1
Xclkbuf_3_2_0_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_144_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21085_ net175 _00854_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20036_ _03275_ _03276_ _05190_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__and3b_1
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _04041_ _04497_ _04518_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__o21ai_4
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ clknet_leaf_1_i_clk _00707_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _04448_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__inv_2
X_20869_ clknet_leaf_93_i_clk _00638_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13410_ _06138_ _06141_ _06146_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__o21a_1
XFILLER_70_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10622_ _03650_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14390_ _07120_ _07126_ vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__xor2_1
XFILLER_139_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13341_ _06045_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__clkbuf_4
XFILLER_195_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10553_ rbzero.tex_r0\[14\] rbzero.tex_r0\[13\] _03613_ vssd1 vssd1 vccd1 vccd1 _03614_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16060_ _07929_ vssd1 vssd1 vccd1 vccd1 _08705_ sky130_fd_sc_hd__buf_4
XFILLER_154_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13272_ _06008_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__clkbuf_4
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _03577_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15011_ _03912_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__clkbuf_4
X_12223_ _04891_ _04992_ _04890_ _04892_ _04969_ _04966_ vssd1 vssd1 vccd1 vccd1 _04993_
+ sky130_fd_sc_hd__mux4_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12154_ _04907_ _04905_ _04921_ _04923_ _04924_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__a2111o_2
XFILLER_162_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ _03903_ vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19750_ _03047_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__clkbuf_4
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12085_ net3 _04852_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__nor2_2
X_16962_ _09470_ _09602_ vssd1 vssd1 vccd1 vccd1 _09603_ sky130_fd_sc_hd__xnor2_1
XFILLER_104_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18701_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.stepDistY\[-12\]
+ _02395_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a21o_1
X_15913_ _08556_ _08552_ vssd1 vssd1 vccd1 vccd1 _08558_ sky130_fd_sc_hd__xor2_1
X_11036_ _03867_ vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__clkbuf_1
X_16893_ _09395_ _09396_ _09397_ _09398_ vssd1 vssd1 vccd1 vccd1 _09534_ sky130_fd_sc_hd__o2bb2a_1
X_19681_ rbzero.pov.spi_buffer\[16\] rbzero.pov.spi_buffer\[17\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03067_ sky130_fd_sc_hd__mux2_1
XFILLER_49_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18632_ _08159_ _09138_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__nor2_1
X_15844_ _08487_ _08488_ vssd1 vssd1 vccd1 vccd1 _08489_ sky130_fd_sc_hd__nand2_1
XFILLER_65_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18563_ _08257_ _09162_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__or2_1
X_15775_ _08054_ _08419_ vssd1 vssd1 vccd1 vccd1 _08420_ sky130_fd_sc_hd__nor2_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _05723_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__inv_2
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ _10070_ _10079_ vssd1 vssd1 vccd1 vccd1 _10080_ sky130_fd_sc_hd__xnor2_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _07462_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__clkbuf_1
X_18494_ _02186_ _02191_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__xor2_1
X_11938_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _04263_ vssd1 vssd1 vccd1 vccd1 _04714_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _09718_ _09720_ vssd1 vssd1 vccd1 vccd1 _10012_ sky130_fd_sc_hd__nor2_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14657_ _07393_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__buf_2
X_11869_ rbzero.tex_g1\[19\] rbzero.tex_g1\[18\] _04336_ vssd1 vssd1 vccd1 vccd1 _04646_
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13608_ _05988_ _06337_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__o21ba_1
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17376_ _09941_ _09942_ vssd1 vssd1 vccd1 vccd1 _09943_ sky130_fd_sc_hd__or2b_1
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14588_ _07116_ _07324_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__or2_1
XFILLER_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16327_ _08180_ _08189_ _08971_ _08170_ vssd1 vssd1 vccd1 vccd1 _08972_ sky130_fd_sc_hd__o22a_1
X_19115_ rbzero.spi_registers.spi_cmd\[0\] rbzero.spi_registers.spi_cmd\[1\] _02690_
+ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__mux2_1
XFILLER_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13539_ _06232_ _06275_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__xor2_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19046_ rbzero.pov.spi_buffer\[54\] rbzero.pov.ready_buffer\[54\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02655_ sky130_fd_sc_hd__mux2_1
X_16258_ _08889_ _08891_ vssd1 vssd1 vccd1 vccd1 _08903_ sky130_fd_sc_hd__nor2_1
XFILLER_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15209_ _07850_ _07854_ _07860_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__and3_1
XFILLER_173_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ _08820_ _08826_ vssd1 vssd1 vccd1 vccd1 _08834_ sky130_fd_sc_hd__nor2_1
XFILLER_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19948_ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__buf_2
XFILLER_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19879_ _03184_ _03187_ _02714_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__o21a_1
XFILLER_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20723_ clknet_leaf_82_i_clk _00492_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_24_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20654_ clknet_leaf_52_i_clk _00438_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_63_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20585_ _07689_ _03454_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__xnor2_1
XFILLER_109_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_78_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21206_ clknet_leaf_26_i_clk _00975_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21137_ clknet_leaf_97_i_clk _00906_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21068_ net158 _00837_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20019_ net59 _03263_ _03264_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__a21oi_1
XFILLER_150_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12910_ _05615_ _05601_ _05566_ _05563_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__o211a_1
XFILLER_207_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13890_ _06626_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__inv_2
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12841_ rbzero.wall_tracer.visualWallDist\[-4\] _05570_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05578_ sky130_fd_sc_hd__a21o_1
XFILLER_74_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_16_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _08194_ _08204_ vssd1 vssd1 vccd1 vccd1 _08205_ sky130_fd_sc_hd__nor2_2
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ rbzero.map_rom.f1 _05517_ _05414_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__mux2_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _07234_ _07246_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__and2_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ gpout0.vpos\[3\] _04041_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__nand2_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _08059_ _08135_ vssd1 vssd1 vccd1 vccd1 _08136_ sky130_fd_sc_hd__nor2_1
XFILLER_42_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.stepDistX\[-12\]
+ _09807_ vssd1 vssd1 vccd1 vccd1 _09809_ sky130_fd_sc_hd__o21ai_1
X_14442_ _07108_ _07063_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__and2b_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11654_ _04422_ _04432_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__nor2_1
XFILLER_122_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ rbzero.tex_g1\[52\] rbzero.tex_g1\[53\] _03635_ vssd1 vssd1 vccd1 vccd1 _03641_
+ sky130_fd_sc_hd__mux2_1
X_17161_ rbzero.traced_texa\[-8\] _09766_ _09767_ rbzero.wall_tracer.visualWallDist\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__a22o_1
XFILLER_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14373_ _07108_ _07109_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__xnor2_2
X_11585_ rbzero.tex_r1\[27\] rbzero.tex_r1\[26\] _04262_ vssd1 vssd1 vccd1 vccd1 _04364_
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16112_ _08725_ _08734_ _08736_ vssd1 vssd1 vccd1 vccd1 _08757_ sky130_fd_sc_hd__and3_1
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13324_ _05944_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__clkbuf_4
XFILLER_70_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10536_ rbzero.tex_r0\[22\] rbzero.tex_r0\[21\] _03602_ vssd1 vssd1 vccd1 vccd1 _03605_
+ sky130_fd_sc_hd__mux2_1
X_17092_ _09476_ _09586_ _09731_ vssd1 vssd1 vccd1 vccd1 _09732_ sky130_fd_sc_hd__a21oi_2
XFILLER_116_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16043_ _08284_ _08128_ _08623_ _08687_ vssd1 vssd1 vccd1 vccd1 _08688_ sky130_fd_sc_hd__o31ai_2
XFILLER_115_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13255_ _05990_ _05991_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__nand2_1
X_10467_ _03568_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__clkbuf_1
X_12206_ net17 _04968_ _04971_ _04975_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__o211a_1
X_13186_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__buf_4
X_10398_ _03530_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__clkbuf_1
X_19802_ rbzero.pov.mosi rbzero.pov.mosi_buffer\[0\] _05189_ vssd1 vssd1 vccd1 vccd1
+ _03130_ sky130_fd_sc_hd__mux2_1
X_12137_ net10 vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__clkinv_2
XFILLER_97_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17994_ _01694_ _01695_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__03302_ clknet_0__03302_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03302_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19733_ _03094_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__clkbuf_1
X_12068_ net2 vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__clkbuf_4
X_16945_ _09583_ _09585_ vssd1 vssd1 vccd1 vccd1 _09586_ sky130_fd_sc_hd__xor2_1
XFILLER_38_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11019_ _03858_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__clkbuf_1
X_19664_ rbzero.pov.spi_buffer\[8\] rbzero.pov.spi_buffer\[9\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03058_ sky130_fd_sc_hd__mux2_1
XFILLER_77_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16876_ _09477_ _09516_ vssd1 vssd1 vccd1 vccd1 _09517_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18615_ _02310_ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__or2_2
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _08471_ _08023_ vssd1 vssd1 vccd1 vccd1 _08472_ sky130_fd_sc_hd__xor2_2
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18546_ _10248_ _01524_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__nor2_1
X_15758_ _08393_ _08395_ vssd1 vssd1 vccd1 vccd1 _08403_ sky130_fd_sc_hd__or2_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ _05742_ _07400_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__nor2_1
X_18477_ _10239_ _09215_ _02173_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__o21ai_1
XFILLER_166_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15689_ _08330_ _08333_ vssd1 vssd1 vccd1 vccd1 _08334_ sky130_fd_sc_hd__nand2_1
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17428_ _05211_ _08215_ _09565_ vssd1 vssd1 vccd1 vccd1 _09995_ sky130_fd_sc_hd__or3_1
XFILLER_178_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17359_ _09924_ _09925_ vssd1 vssd1 vccd1 vccd1 _09926_ sky130_fd_sc_hd__xnor2_1
XFILLER_158_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19029_ rbzero.pov.spi_buffer\[46\] rbzero.pov.ready_buffer\[46\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02646_ sky130_fd_sc_hd__mux2_1
XFILLER_173_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20114__147 clknet_1_1__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__inv_2
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20706_ clknet_leaf_51_i_clk _00490_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20195__219 clknet_1_1__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__inv_2
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20637_ clknet_leaf_65_i_clk _00421_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11370_ rbzero.row_render.size\[3\] _04149_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__or2_1
XFILLER_166_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20568_ rbzero.traced_texVinit\[11\] _03443_ _07756_ _01552_ vssd1 vssd1 vccd1 vccd1
+ _01419_ sky130_fd_sc_hd__a22o_1
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10321_ rbzero.tex_r1\[57\] rbzero.tex_r1\[58\] _03483_ vssd1 vssd1 vccd1 vccd1 _03490_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20499_ _03390_ _03394_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__nand2_1
X_13040_ _05776_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__clkbuf_2
XFILLER_106_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20089__124 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__inv_2
XFILLER_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14991_ rbzero.wall_tracer.stepDistX\[2\] _07562_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07666_ sky130_fd_sc_hd__mux2_1
XFILLER_94_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16730_ _09363_ _09371_ vssd1 vssd1 vccd1 vccd1 _09372_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13942_ _06675_ _06678_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__nor2_1
XFILLER_120_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16661_ _09299_ _09300_ _09302_ vssd1 vssd1 vccd1 vccd1 _09304_ sky130_fd_sc_hd__a21o_1
X_13873_ _06609_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18400_ _02083_ _02098_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__xnor2_1
X_15612_ _08214_ vssd1 vssd1 vccd1 vccd1 _08257_ sky130_fd_sc_hd__clkbuf_4
X_12824_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__clkbuf_4
X_16592_ _09231_ _09233_ vssd1 vssd1 vccd1 vccd1 _09235_ sky130_fd_sc_hd__and2_1
X_19380_ rbzero.wall_tracer.rayAddendY\[-2\] _00013_ _02867_ vssd1 vssd1 vccd1 vccd1
+ _00808_ sky130_fd_sc_hd__o21a_1
XFILLER_163_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18331_ _01646_ _01972_ _10271_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a21o_1
X_15543_ _08148_ _08183_ _08185_ _08187_ vssd1 vssd1 vccd1 vccd1 _08188_ sky130_fd_sc_hd__a31o_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12755_ _05502_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__clkbuf_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18262_ _01839_ _01847_ _01961_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__a21oi_2
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ rbzero.debug_overlay.facingY\[-5\] _04454_ _04463_ rbzero.debug_overlay.facingY\[-3\]
+ _04484_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__a221o_1
XFILLER_202_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15474_ _08064_ _08118_ vssd1 vssd1 vccd1 vccd1 _08119_ sky130_fd_sc_hd__xnor2_1
XFILLER_124_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12686_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__or2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14425_ _07144_ _07161_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__nand2_1
X_17213_ _09791_ _09794_ vssd1 vssd1 vccd1 vccd1 _09795_ sky130_fd_sc_hd__xnor2_1
X_18193_ _01892_ _01893_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__nand2_1
XFILLER_202_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11637_ gpout0.hpos\[3\] _04023_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__nor2_1
XFILLER_129_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17144_ _07549_ _09763_ rbzero.row_render.size\[6\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00534_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_129_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14356_ _07090_ _07092_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__nor2_1
XFILLER_156_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11568_ _04135_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__buf_4
XFILLER_7_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ _06040_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10519_ rbzero.tex_r0\[30\] rbzero.tex_r0\[29\] _03591_ vssd1 vssd1 vccd1 vccd1 _03596_
+ sky130_fd_sc_hd__mux2_1
X_17075_ _09567_ _09569_ vssd1 vssd1 vccd1 vccd1 _09715_ sky130_fd_sc_hd__nor2_1
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14287_ _06784_ _06796_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__or2b_1
X_11499_ rbzero.tex_r0\[13\] rbzero.tex_r0\[12\] _04273_ vssd1 vssd1 vccd1 vccd1 _04279_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16026_ _08620_ _08670_ vssd1 vssd1 vccd1 vccd1 _08671_ sky130_fd_sc_hd__nor2_1
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13238_ _05889_ _05899_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__xnor2_4
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13169_ _05863_ _05868_ _05811_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__mux2_1
XFILLER_151_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17977_ _01555_ _01557_ _01554_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__a21boi_2
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19716_ _03085_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_66_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16928_ _09428_ _09435_ _09568_ vssd1 vssd1 vccd1 vccd1 _09569_ sky130_fd_sc_hd__a21oi_2
XFILLER_133_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03316_ _03316_ vssd1 vssd1 vccd1 vccd1 clknet_0__03316_ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19647_ _03049_ vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16859_ _09387_ _09390_ vssd1 vssd1 vccd1 vccd1 _09500_ sky130_fd_sc_hd__nand2_1
XFILLER_20_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18529_ _02125_ _02128_ _02225_ _05203_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__a31o_1
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21540_ net461 _01309_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21471_ net392 _01240_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20422_ _09750_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__clkbuf_4
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10870_ _03780_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__and2_1
XFILLER_101_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ _05223_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__and2b_1
Xclkbuf_1_0__f__03305_ clknet_0__03305_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03305_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14210_ _06664_ _06940_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__nand2_1
X_11422_ _04175_ _04177_ _04201_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _04202_
+ sky130_fd_sc_hd__o2bb2a_1
X_15190_ _07820_ rbzero.wall_tracer.rayAddendX\[7\] vssd1 vssd1 vccd1 vccd1 _07843_
+ sky130_fd_sc_hd__nand2_1
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14141_ _06858_ _06876_ _06877_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__a21boi_1
X_11353_ rbzero.floor_leak\[3\] _04119_ _04121_ rbzero.floor_leak\[4\] _04132_ vssd1
+ vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__a221o_1
XFILLER_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ net45 net44 vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__xor2_4
XFILLER_153_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14072_ _06806_ _06808_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__nand2_1
XFILLER_141_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11284_ _04062_ _04061_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__nand2_1
XFILLER_193_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17900_ _01472_ _01484_ _01482_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__a21oi_1
X_13023_ _05695_ _05702_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__or2_1
XFILLER_112_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18880_ _02550_ _02551_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17831_ _01513_ _01534_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__xnor2_2
XFILLER_121_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17762_ _01464_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__xnor2_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14974_ rbzero.wall_tracer.stepDistX\[-6\] _07650_ vssd1 vssd1 vccd1 vccd1 _07657_
+ sky130_fd_sc_hd__nor2_1
XFILLER_94_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19501_ _02905_ rbzero.debug_overlay.vplaneY\[-1\] vssd1 vssd1 vccd1 vccd1 _02980_
+ sky130_fd_sc_hd__or2_1
XFILLER_207_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16713_ _08054_ _09164_ vssd1 vssd1 vccd1 vccd1 _09355_ sky130_fd_sc_hd__nor2_1
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13925_ _06661_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__clkbuf_2
X_17693_ _10137_ _10141_ _10140_ vssd1 vssd1 vccd1 vccd1 _10258_ sky130_fd_sc_hd__a21bo_1
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19432_ _02899_ _02915_ _02914_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a21o_1
X_16644_ _05194_ _09285_ _09286_ _08224_ vssd1 vssd1 vccd1 vccd1 _09287_ sky130_fd_sc_hd__a31o_1
X_13856_ _06567_ _06592_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12807_ _05533_ _05546_ _05547_ _05284_ rbzero.wall_tracer.mapY\[8\] vssd1 vssd1
+ vccd1 vccd1 _00415_ sky130_fd_sc_hd__a32o_1
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19363_ _04471_ rbzero.wall_tracer.rayAddendY\[-3\] vssd1 vssd1 vccd1 vccd1 _02852_
+ sky130_fd_sc_hd__nand2_1
XFILLER_188_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16575_ _08162_ _09217_ vssd1 vssd1 vccd1 vccd1 _09218_ sky130_fd_sc_hd__nor2_1
X_13787_ _06507_ _06523_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__nor2_1
XFILLER_188_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10999_ rbzero.tex_b0\[58\] rbzero.tex_b0\[57\] _03843_ vssd1 vssd1 vccd1 vccd1 _03848_
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20143__173 clknet_1_0__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__inv_2
XFILLER_16_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18314_ _01903_ _01906_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__nor2_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _05434_ _05485_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__nand2_1
X_15526_ _07549_ _07552_ _07555_ vssd1 vssd1 vccd1 vccd1 _08171_ sky130_fd_sc_hd__a21oi_4
XFILLER_203_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19294_ rbzero.spi_registers.new_other\[1\] rbzero.spi_registers.spi_buffer\[1\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__mux2_1
XFILLER_188_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18245_ _09661_ _09359_ _01829_ _01944_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__o31a_1
X_15457_ _07925_ _08100_ _08101_ vssd1 vssd1 vccd1 vccd1 _08102_ sky130_fd_sc_hd__a21oi_4
X_12669_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__or2_1
XFILLER_198_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14408_ _06680_ _06761_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__nor2_1
XFILLER_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18176_ _01758_ _01760_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__nand2_1
XFILLER_128_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15388_ _07990_ _08032_ vssd1 vssd1 vccd1 vccd1 _08033_ sky130_fd_sc_hd__nand2_1
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17127_ _04154_ _04442_ vssd1 vssd1 vccd1 vccd1 _09758_ sky130_fd_sc_hd__or2_1
XFILLER_143_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14339_ _07071_ _07074_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__or2_1
XFILLER_116_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17058_ _07585_ _09697_ _09431_ _09085_ vssd1 vssd1 vccd1 vccd1 _09698_ sky130_fd_sc_hd__a31o_1
XFILLER_143_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16009_ _08622_ _08653_ vssd1 vssd1 vccd1 vccd1 _08654_ sky130_fd_sc_hd__xor2_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20971_ clknet_leaf_12_i_clk _00740_ vssd1 vssd1 vccd1 vccd1 rbzero.floor_leak\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20226__248 clknet_1_0__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__inv_2
XFILLER_199_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21523_ net444 _01292_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21454_ net375 _01223_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21385_ net306 _01154_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput58 net58 vssd1 vssd1 vccd1 vccd1 o_gpout[5] sky130_fd_sc_hd__clkbuf_1
Xoutput69 net69 vssd1 vssd1 vccd1 vccd1 o_tex_out0 sky130_fd_sc_hd__buf_2
XFILLER_27_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11971_ rbzero.tex_b1\[27\] rbzero.tex_b1\[26\] _04262_ vssd1 vssd1 vccd1 vccd1 _04746_
+ sky130_fd_sc_hd__mux2_1
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _06078_ _06016_ _06445_ _06446_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__o31a_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10922_ rbzero.tex_b1\[30\] rbzero.tex_b1\[31\] _03806_ vssd1 vssd1 vccd1 vccd1 _03808_
+ sky130_fd_sc_hd__mux2_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _07343_ _07344_ _07346_ _07378_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__o211ai_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ _06279_ _06377_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__nand2_1
XFILLER_72_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10853_ _03771_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _09003_ _09004_ vssd1 vssd1 vccd1 vccd1 _09005_ sky130_fd_sc_hd__nand2_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13572_ _06103_ _06104_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__xnor2_1
X_10784_ _03735_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _07951_ _07955_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__nand2_1
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _05213_ _05232_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__o21a_4
X_16291_ _08911_ _08934_ _08935_ vssd1 vssd1 vccd1 vccd1 _08936_ sky130_fd_sc_hd__o21ba_1
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18030_ _01700_ _01731_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__xor2_1
X_15242_ _04035_ _07889_ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__and2_1
XFILLER_173_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12454_ _05208_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__clkbuf_4
XFILLER_185_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11405_ rbzero.row_render.size\[4\] _04150_ rbzero.row_render.size\[5\] vssd1 vssd1
+ vccd1 vccd1 _04185_ sky130_fd_sc_hd__o21ai_1
XFILLER_158_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15173_ _07827_ vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__clkbuf_1
X_12385_ _05145_ _05146_ gpout5.clk_div\[1\] _05151_ net34 vssd1 vssd1 vccd1 vccd1
+ _05152_ sky130_fd_sc_hd__a311o_2
XFILLER_193_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14124_ _06825_ _06832_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__xnor2_1
XFILLER_197_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11336_ _04114_ _04115_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__or2_4
X_19981_ rbzero.pov.ready_buffer\[30\] _03252_ _03253_ rbzero.debug_overlay.facingY\[-1\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__o221a_1
X_20173__199 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__inv_2
XFILLER_125_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14055_ _06778_ _06790_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__nand2_1
X_18932_ _02594_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__clkbuf_4
X_11267_ gpout0.vpos\[6\] _04043_ _04044_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_
+ sky130_fd_sc_hd__a211o_4
XFILLER_158_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13006_ _05700_ _05732_ _05738_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__nor3b_2
XFILLER_80_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18863_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.stepDistY\[9\] vssd1
+ vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__or2_1
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11198_ _03972_ _03980_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__or3b_4
XFILLER_95_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17814_ _09434_ _09988_ _08895_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__a21oi_1
XFILLER_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18794_ rbzero.wall_tracer.trackDistY\[-1\] _02477_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02478_ sky130_fd_sc_hd__mux2_1
XFILLER_48_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17745_ _01445_ _01447_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__or2_1
XFILLER_36_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14957_ rbzero.wall_tracer.visualWallDist\[10\] _07594_ vssd1 vssd1 vccd1 vccd1 _07648_
+ sky130_fd_sc_hd__or2_1
X_13908_ _06574_ _06585_ _06634_ _06635_ _06636_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__a32o_1
X_17676_ _10237_ _10240_ vssd1 vssd1 vccd1 vccd1 _10241_ sky130_fd_sc_hd__nand2_1
X_14888_ _07591_ _07597_ _07599_ _04039_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__o211a_1
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19415_ _02887_ _02890_ _02898_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__nand3_1
X_16627_ _08283_ _08189_ vssd1 vssd1 vccd1 vccd1 _09270_ sky130_fd_sc_hd__nor2_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13839_ _06015_ _05991_ _05978_ _06055_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__or4_1
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19346_ _02827_ _02835_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a21boi_1
X_16558_ _09082_ _09201_ vssd1 vssd1 vccd1 vccd1 _09202_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15509_ _08152_ _08153_ vssd1 vssd1 vccd1 vccd1 _08154_ sky130_fd_sc_hd__or2_1
XFILLER_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19277_ _02793_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16489_ _07602_ _08230_ _08147_ _08236_ vssd1 vssd1 vccd1 vccd1 _09133_ sky130_fd_sc_hd__or4_1
XFILLER_50_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18228_ _01811_ _01927_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18159_ _08237_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__clkbuf_4
XFILLER_172_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21170_ clknet_leaf_92_i_clk _00939_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20052_ _04890_ _04037_ _03287_ _03911_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__a31o_1
XFILLER_131_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20954_ clknet_leaf_94_i_clk _00723_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20885_ clknet_leaf_88_i_clk _00654_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21506_ net427 _01275_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21437_ net358 _01206_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12170_ net42 _04918_ _04905_ _04940_ net12 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__a311o_1
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21368_ net289 _01137_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11121_ _03555_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__buf_6
XFILLER_162_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21299_ net220 _01068_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11052_ _03875_ vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _08492_ _08494_ _08503_ _08504_ vssd1 vssd1 vccd1 vccd1 _08505_ sky130_fd_sc_hd__a31o_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14811_ _07459_ _07404_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__nor2_1
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20209__232 clknet_1_0__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__inv_2
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _08406_ _08414_ _08434_ vssd1 vssd1 vccd1 vccd1 _08436_ sky130_fd_sc_hd__nand3_1
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _10093_ _10095_ vssd1 vssd1 vccd1 vccd1 _10096_ sky130_fd_sc_hd__nand2_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20361__369 clknet_1_0__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__inv_2
X_14742_ _05807_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__clkbuf_4
X_11954_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _04356_ vssd1 vssd1 vccd1 vccd1 _04730_
+ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_104 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_104/HI zeros[14]
+ sky130_fd_sc_hd__conb_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_115 vssd1 vssd1 vccd1 vccd1 ones[9] top_ew_algofoogle_115/LO sky130_fd_sc_hd__conb_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10905_ rbzero.tex_b1\[38\] rbzero.tex_b1\[39\] _03795_ vssd1 vssd1 vccd1 vccd1 _03799_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14673_ _07409_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__inv_2
X_17461_ _09889_ _10027_ vssd1 vssd1 vccd1 vccd1 _10028_ sky130_fd_sc_hd__or2_1
X_11885_ _04140_ _04645_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__or3_1
XFILLER_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19200_ _09753_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__and2_1
X_16412_ _08439_ _08468_ vssd1 vssd1 vccd1 vccd1 _09057_ sky130_fd_sc_hd__nor2_1
X_13624_ _05846_ _05975_ _06285_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__or3_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10836_ rbzero.tex_g0\[8\] rbzero.tex_g0\[7\] _03762_ vssd1 vssd1 vccd1 vccd1 _03763_
+ sky130_fd_sc_hd__mux2_1
X_17392_ _08445_ _08332_ vssd1 vssd1 vccd1 vccd1 _09959_ sky130_fd_sc_hd__nand2_1
XFILLER_60_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19131_ _02700_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__clkbuf_1
XFILLER_164_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16343_ _08977_ _08243_ vssd1 vssd1 vccd1 vccd1 _08988_ sky130_fd_sc_hd__or2_1
X_13555_ _05995_ _06113_ _06061_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__a21o_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10767_ _03726_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ _05255_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.trackDistX\[0\]
+ _05257_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__a22o_1
XFILLER_201_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16274_ _08915_ _08918_ vssd1 vssd1 vccd1 vccd1 _08919_ sky130_fd_sc_hd__xor2_1
XFILLER_121_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19062_ _02663_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__clkbuf_1
X_13486_ _06183_ _06222_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__xor2_1
X_10698_ rbzero.tex_g1\[8\] rbzero.tex_g1\[9\] _03680_ vssd1 vssd1 vccd1 vccd1 _03690_
+ sky130_fd_sc_hd__mux2_1
XFILLER_172_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18013_ _01705_ _01714_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__xor2_1
X_15225_ _07742_ _07730_ _07862_ _07821_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__a211oi_1
XFILLER_173_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12437_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__clkinv_4
X_20255__274 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__inv_2
XFILLER_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15156_ _07811_ vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__clkbuf_1
X_12368_ _05121_ _05135_ net31 vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__and3b_1
XFILLER_126_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14107_ _05825_ _06668_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__nor2_1
XFILLER_10_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11319_ _04098_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__inv_2
X_15087_ _07741_ _07745_ _07746_ vssd1 vssd1 vccd1 vccd1 _07747_ sky130_fd_sc_hd__a21oi_1
X_19964_ rbzero.pov.ready_buffer\[38\] _03247_ _03249_ rbzero.debug_overlay.facingX\[-4\]
+ _03250_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__a221o_1
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12299_ _05044_ _05047_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__nand2_1
XFILLER_141_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18915_ _02582_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__clkbuf_1
X_14038_ _06771_ _06772_ _06773_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__o21bai_1
XFILLER_171_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19895_ rbzero.debug_overlay.playerY\[-8\] _03198_ _03200_ _03157_ vssd1 vssd1 vccd1
+ vccd1 _00990_ sky130_fd_sc_hd__o211a_1
XFILLER_84_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18846_ rbzero.wall_tracer.trackDistY\[6\] _02522_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02523_ sky130_fd_sc_hd__mux2_1
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18777_ rbzero.wall_tracer.trackDistY\[-3\] _02462_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02463_ sky130_fd_sc_hd__mux2_1
XFILLER_110_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15989_ _08630_ _08631_ _08632_ _08633_ vssd1 vssd1 vccd1 vccd1 _08634_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17728_ _10289_ _10291_ vssd1 vssd1 vccd1 vccd1 _10293_ sky130_fd_sc_hd__and2_1
XFILLER_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17659_ _10222_ _10223_ vssd1 vssd1 vccd1 vccd1 _10224_ sky130_fd_sc_hd__and2b_1
XFILLER_63_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20670_ clknet_leaf_61_i_clk _00454_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_195_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19329_ _02728_ _02820_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__or2_1
XFILLER_104_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21222_ clknet_leaf_21_i_clk _00991_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21153_ clknet_leaf_87_i_clk _00922_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21084_ net174 _00853_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20035_ _04021_ _04026_ _02705_ _04989_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__a31o_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20937_ clknet_leaf_93_i_clk _00706_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11670_ _04427_ _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__nor2_1
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20868_ clknet_leaf_5_i_clk _00637_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10621_ rbzero.tex_g1\[45\] rbzero.tex_g1\[46\] _03647_ vssd1 vssd1 vccd1 vccd1 _03650_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20799_ clknet_leaf_44_i_clk _00568_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13340_ _06040_ _06043_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__a21oi_1
X_10552_ _03557_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13271_ _05946_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__or2_1
X_10483_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _03569_ vssd1 vssd1 vccd1 vccd1 _03577_
+ sky130_fd_sc_hd__mux2_1
X_15010_ _07675_ vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12222_ gpout0.vpos\[0\] vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__buf_2
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12153_ clknet_1_1__leaf__04835_ _04918_ _04905_ vssd1 vssd1 vccd1 vccd1 _04924_
+ sky130_fd_sc_hd__and3_2
XFILLER_151_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ rbzero.tex_b0\[8\] rbzero.tex_b0\[7\] _03898_ vssd1 vssd1 vccd1 vccd1 _03903_
+ sky130_fd_sc_hd__mux2_1
XFILLER_190_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12084_ net46 _04853_ _04854_ _04855_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__a22o_1
X_16961_ _09082_ _09601_ vssd1 vssd1 vccd1 vccd1 _09602_ sky130_fd_sc_hd__xnor2_1
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18700_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.stepDistY\[-12\]
+ _09807_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__o21ai_1
X_15912_ _08552_ _08556_ vssd1 vssd1 vccd1 vccd1 _08557_ sky130_fd_sc_hd__or2b_1
X_11035_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _03865_ vssd1 vssd1 vccd1 vccd1 _03867_
+ sky130_fd_sc_hd__mux2_1
X_19680_ _03066_ vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__clkbuf_1
X_16892_ _09531_ _09532_ vssd1 vssd1 vccd1 vccd1 _09533_ sky130_fd_sc_hd__xnor2_2
XFILLER_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18631_ _02271_ _02280_ _02278_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a21oi_1
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _08478_ _08485_ _08486_ vssd1 vssd1 vccd1 vccd1 _08488_ sky130_fd_sc_hd__nand3_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18562_ _02257_ _02258_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__xnor2_2
XFILLER_92_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _08417_ _08418_ vssd1 vssd1 vccd1 vccd1 _08419_ sky130_fd_sc_hd__nand2_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _05670_ _05671_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__nand2_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _10072_ _10078_ vssd1 vssd1 vccd1 vccd1 _10079_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14725_ rbzero.wall_tracer.stepDistY\[-12\] _07460_ _07461_ vssd1 vssd1 vccd1 vccd1
+ _07462_ sky130_fd_sc_hd__mux2_1
XFILLER_205_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18493_ _02189_ _02190_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__xor2_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ rbzero.tex_b0\[55\] _04221_ _04222_ _04218_ vssd1 vssd1 vccd1 vccd1 _04713_
+ sky130_fd_sc_hd__a31o_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _09972_ _10010_ vssd1 vssd1 vccd1 vccd1 _10011_ sky130_fd_sc_hd__xnor2_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11868_ _04371_ _04632_ _04636_ _04644_ _04244_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__o311a_1
X_14656_ _05703_ _05928_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__or2_1
XFILLER_20_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13607_ _06338_ _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__and2b_1
XFILLER_32_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10819_ rbzero.tex_g0\[16\] rbzero.tex_g0\[15\] _03751_ vssd1 vssd1 vccd1 vccd1 _03754_
+ sky130_fd_sc_hd__mux2_1
X_17375_ _09522_ _08705_ _08419_ vssd1 vssd1 vccd1 vccd1 _09942_ sky130_fd_sc_hd__or3_1
X_11799_ rbzero.tex_g0\[46\] _04336_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__and2_1
X_14587_ _06696_ _07072_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__and2_1
XFILLER_159_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19114_ _02691_ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16326_ _05209_ rbzero.wall_tracer.stepDistX\[3\] _08214_ vssd1 vssd1 vccd1 vccd1
+ _08971_ sky130_fd_sc_hd__a21boi_2
XFILLER_159_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13538_ _06273_ _06274_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__nor2_1
XFILLER_185_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19045_ _02654_ vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16257_ _08836_ _08842_ vssd1 vssd1 vccd1 vccd1 _08902_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13469_ _06154_ _06205_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15208_ _07742_ _07847_ _07859_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__a21o_1
XFILLER_12_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16188_ _08828_ _08832_ vssd1 vssd1 vccd1 vccd1 _08833_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15139_ rbzero.wall_tracer.rayAddendX\[3\] _07695_ _07795_ _07703_ vssd1 vssd1 vccd1
+ vccd1 _07796_ sky130_fd_sc_hd__a22o_1
XFILLER_5_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19947_ rbzero.pov.ready _02708_ _02820_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__nand3_4
XFILLER_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19878_ rbzero.pov.ready_buffer\[72\] _03164_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_
+ sky130_fd_sc_hd__o21a_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18829_ _09863_ _02506_ _02507_ _01677_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__o31ai_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20722_ clknet_leaf_80_i_clk _00491_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20653_ clknet_leaf_56_i_clk _00437_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20584_ _07684_ _07690_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__and2b_1
XFILLER_20_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21205_ clknet_leaf_23_i_clk _00974_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21136_ clknet_leaf_97_i_clk _00905_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21067_ net157 _00836_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20018_ _04006_ _04811_ _04813_ _03262_ _03911_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a41o_1
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12840_ _05561_ _05468_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__or2_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ rbzero.debug_overlay.playerX\[3\] _05516_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05517_ sky130_fd_sc_hd__mux2_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _07234_ _07246_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__nor2_1
X_11722_ rbzero.debug_overlay.playerY\[2\] _04451_ _04466_ rbzero.debug_overlay.playerY\[-8\]
+ _04500_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__a221o_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19573__30 clknet_1_1__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__inv_2
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _07951_ _08133_ _08134_ _05197_ vssd1 vssd1 vccd1 vccd1 _08135_ sky130_fd_sc_hd__o211ai_4
XFILLER_199_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _07109_ _07177_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11653_ _04430_ _04431_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__or2b_1
XFILLER_187_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10604_ _03640_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14372_ _06240_ _06658_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__or2_1
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17160_ rbzero.traced_texa\[-9\] _09766_ _09767_ rbzero.wall_tracer.visualWallDist\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__a22o_1
X_11584_ _04359_ _04362_ _04332_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__mux2_1
XFILLER_122_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16111_ _08740_ _08755_ vssd1 vssd1 vccd1 vccd1 _08756_ sky130_fd_sc_hd__nand2_1
X_13323_ _05923_ _05989_ _05983_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__a21bo_1
XFILLER_196_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10535_ _03604_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__clkbuf_1
X_17091_ _09583_ _09585_ vssd1 vssd1 vccd1 vccd1 _09731_ sky130_fd_sc_hd__nor2_1
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16042_ _08684_ _08686_ vssd1 vssd1 vccd1 vccd1 _08687_ sky130_fd_sc_hd__or2b_1
X_13254_ _05920_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10466_ rbzero.tex_r0\[55\] rbzero.tex_r0\[54\] _03558_ vssd1 vssd1 vccd1 vccd1 _03568_
+ sky130_fd_sc_hd__mux2_1
XFILLER_129_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12205_ _04960_ net16 _04972_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__and4_1
X_13185_ _05889_ _05900_ _05910_ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a31o_1
X_10397_ rbzero.tex_r1\[21\] rbzero.tex_r1\[22\] _03527_ vssd1 vssd1 vccd1 vccd1 _03530_
+ sky130_fd_sc_hd__mux2_1
X_19801_ _03129_ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__clkbuf_1
X_12136_ _04906_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__buf_4
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17993_ _01687_ _01609_ _01693_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__and3_1
XFILLER_111_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03301_ clknet_0__03301_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03301_
+ sky130_fd_sc_hd__clkbuf_16
X_19732_ rbzero.pov.spi_buffer\[40\] rbzero.pov.spi_buffer\[41\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03094_ sky130_fd_sc_hd__mux2_1
X_12067_ _04837_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nand2_1
X_16944_ _09382_ _09447_ _09584_ vssd1 vssd1 vccd1 vccd1 _09585_ sky130_fd_sc_hd__a21oi_1
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20367__375 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__inv_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11018_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _03854_ vssd1 vssd1 vccd1 vccd1 _03858_
+ sky130_fd_sc_hd__mux2_1
X_19663_ _03057_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__clkbuf_1
X_16875_ _09514_ _09515_ vssd1 vssd1 vccd1 vccd1 _09516_ sky130_fd_sc_hd__nand2_1
XFILLER_38_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20066__103 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__inv_2
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18614_ _02307_ _02309_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__and2_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _08024_ _08014_ vssd1 vssd1 vccd1 vccd1 _08471_ sky130_fd_sc_hd__nand2_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18545_ _10248_ _10266_ _02151_ _02045_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__o31a_1
X_15757_ _08064_ _08118_ _08401_ vssd1 vssd1 vccd1 vccd1 _08402_ sky130_fd_sc_hd__a21o_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _05563_ _05566_ _05591_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__and3_1
XFILLER_79_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14708_ _05779_ _07428_ _07429_ _05742_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__o211a_1
X_18476_ _10239_ _09215_ _02173_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__or3_1
XFILLER_127_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15688_ _08129_ _08104_ _08331_ _08332_ vssd1 vssd1 vccd1 vccd1 _08333_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17427_ _09987_ _09993_ vssd1 vssd1 vccd1 vccd1 _09994_ sky130_fd_sc_hd__xor2_2
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14639_ _05742_ _05755_ _07105_ _07374_ _07375_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__a32o_1
XFILLER_159_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17358_ _08416_ _09704_ vssd1 vssd1 vccd1 vccd1 _09925_ sky130_fd_sc_hd__nor2_1
XFILLER_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16309_ _08619_ _08950_ _08946_ vssd1 vssd1 vccd1 vccd1 _08954_ sky130_fd_sc_hd__and3b_1
XFILLER_173_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ rbzero.wall_tracer.trackDistX\[-6\] _09861_ _05413_ vssd1 vssd1 vccd1 vccd1
+ _09862_ sky130_fd_sc_hd__mux2_1
XFILLER_162_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19028_ _02645_ vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__clkbuf_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20705_ clknet_leaf_56_i_clk _00489_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_200_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03321_ clknet_0__03321_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03321_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20636_ clknet_leaf_64_i_clk _00420_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20567_ rbzero.traced_texVinit\[10\] _03443_ _09771_ _10297_ vssd1 vssd1 vccd1 vccd1
+ _01418_ sky130_fd_sc_hd__a22o_1
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10320_ _03489_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20498_ rbzero.traced_texa\[2\] rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 _03396_
+ sky130_fd_sc_hd__nand2_1
XFILLER_124_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21119_ net209 _00888_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[59\] sky130_fd_sc_hd__dfxtp_1
X_19625__78 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__inv_2
X_14990_ _07665_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_59_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13941_ _06677_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__clkbuf_4
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16660_ _09299_ _09300_ _09302_ vssd1 vssd1 vccd1 vccd1 _09303_ sky130_fd_sc_hd__nand3_1
XFILLER_207_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13872_ _06548_ _06608_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__or2_1
XFILLER_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15611_ _08253_ _08255_ vssd1 vssd1 vccd1 vccd1 _08256_ sky130_fd_sc_hd__xnor2_1
X_12823_ rbzero.wall_tracer.rcp_sel\[0\] vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__clkinv_2
X_16591_ _09231_ _09233_ vssd1 vssd1 vccd1 vccd1 _09234_ sky130_fd_sc_hd__nor2_1
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18330_ _01646_ _02028_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _07951_ _08186_ _05207_ vssd1 vssd1 vccd1 vccd1 _08187_ sky130_fd_sc_hd__a21o_1
XFILLER_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12754_ rbzero.map_rom.f3 _05501_ _05414_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__mux2_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18261_ _01846_ _01840_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__and2b_1
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11705_ rbzero.debug_overlay.facingY\[0\] _04459_ _04460_ rbzero.debug_overlay.facingY\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__a22o_1
XFILLER_91_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15473_ _08108_ _08117_ vssd1 vssd1 vccd1 vccd1 _08118_ sky130_fd_sc_hd__xor2_1
X_12685_ _05431_ _05432_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__and2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17212_ _09792_ _09793_ vssd1 vssd1 vccd1 vccd1 _09794_ sky130_fd_sc_hd__or2_1
X_11636_ gpout0.hpos\[9\] _04414_ _04046_ _04020_ vssd1 vssd1 vccd1 vccd1 _04415_
+ sky130_fd_sc_hd__a211o_2
X_14424_ _07133_ _07143_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__nand2_1
X_18192_ _01890_ _01891_ _01855_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__a21o_1
XFILLER_175_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17143_ _09765_ _09763_ rbzero.row_render.size\[5\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00533_ sky130_fd_sc_hd__a2bb2o_1
X_11567_ _04343_ _04344_ _04345_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__mux2_1
XFILLER_129_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14355_ _06735_ _07030_ _07091_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10518_ _03595_ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__clkbuf_1
X_13306_ _05943_ _06042_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__and2_1
X_17074_ _09702_ _09713_ vssd1 vssd1 vccd1 vccd1 _09714_ sky130_fd_sc_hd__xnor2_4
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14286_ _07015_ _07022_ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__xnor2_2
XFILLER_115_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11498_ rbzero.tex_r0\[15\] _04221_ _04222_ _04219_ vssd1 vssd1 vccd1 vccd1 _04278_
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13237_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__buf_2
X_16025_ _08666_ _08668_ _08669_ vssd1 vssd1 vccd1 vccd1 _08670_ sky130_fd_sc_hd__o21a_1
X_10449_ _03559_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13168_ _05902_ _05874_ _05904_ _05755_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__o22a_1
XFILLER_112_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12119_ gpout0.vpos\[8\] vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__buf_2
XFILLER_97_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13099_ _05640_ _05648_ _05791_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__mux2_1
X_17976_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] vssd1
+ vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__and2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19715_ rbzero.pov.spi_buffer\[32\] rbzero.pov.spi_buffer\[33\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03085_ sky130_fd_sc_hd__mux2_1
X_16927_ _08215_ _09294_ _09427_ vssd1 vssd1 vccd1 vccd1 _09568_ sky130_fd_sc_hd__nor3_1
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_62_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03315_ _03315_ vssd1 vssd1 vccd1 vccd1 clknet_0__03315_ sky130_fd_sc_hd__clkbuf_16
X_19646_ rbzero.pov.mosi rbzero.pov.spi_buffer\[0\] _03048_ vssd1 vssd1 vccd1 vccd1
+ _03049_ sky130_fd_sc_hd__mux2_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16858_ _09366_ _09369_ _09365_ vssd1 vssd1 vccd1 vccd1 _09499_ sky130_fd_sc_hd__a21bo_1
X_20395__20 clknet_1_1__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__inv_2
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15809_ _08444_ _08450_ vssd1 vssd1 vccd1 vccd1 _08454_ sky130_fd_sc_hd__nor2_1
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16789_ _07575_ _08983_ _09430_ vssd1 vssd1 vccd1 vccd1 _09431_ sky130_fd_sc_hd__nor3_2
XFILLER_18_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_77_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18528_ _02125_ _02128_ _02225_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18459_ _02155_ _02156_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__nor2_1
XFILLER_194_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21470_ net391 _01239_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[49\] sky130_fd_sc_hd__dfxtp_1
X_20120__152 clknet_1_0__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__inv_2
XFILLER_21_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20421_ _03272_ _03330_ _03331_ _03327_ rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1
+ _01385_ sky130_fd_sc_hd__a32o_1
XFILLER_101_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_15_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20283_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__buf_1
XFILLER_136_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20203__227 clknet_1_1__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__inv_2
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12470_ rbzero.wall_tracer.trackDistY\[5\] _05222_ _05224_ rbzero.wall_tracer.trackDistY\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__o22ai_1
XFILLER_197_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21668_ clknet_leaf_34_i_clk _01437_ vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__03304_ clknet_0__03304_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03304_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11421_ _04154_ _04179_ _04180_ _04181_ _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__o221a_1
XFILLER_71_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20619_ clknet_leaf_15_i_clk _00403_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.b6 sky130_fd_sc_hd__dfxtp_1
XFILLER_137_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21599_ net140 _01368_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[50\] sky130_fd_sc_hd__dfxtp_1
X_14140_ _06859_ _06875_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__or2b_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11352_ rbzero.floor_leak\[2\] _04123_ _04119_ rbzero.floor_leak\[3\] _04131_ vssd1
+ vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__o221a_1
XFILLER_67_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10303_ _03476_ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__and2_1
X_14071_ _06776_ _06739_ _06804_ _06807_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__o31a_1
X_11283_ rbzero.texV\[6\] _04061_ _04062_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__a21boi_1
XFILLER_141_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13022_ _05756_ _05758_ _05737_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__a21oi_1
XFILLER_79_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17830_ _01532_ _01533_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__and2b_1
XFILLER_126_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17761_ _09391_ _09359_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__nor2_1
X_14973_ _00008_ _07524_ _07656_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__a21oi_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19500_ _02952_ _02976_ _02977_ _02975_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a31o_1
X_16712_ _08331_ _09353_ vssd1 vssd1 vccd1 vccd1 _09354_ sky130_fd_sc_hd__nand2_1
X_13924_ _06613_ _06660_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__or2_1
X_17692_ _09974_ _10255_ _10256_ _10117_ vssd1 vssd1 vccd1 vccd1 _10257_ sky130_fd_sc_hd__a22o_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19431_ _02890_ _02898_ _02885_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a21bo_1
X_16643_ _07575_ _07579_ _08983_ vssd1 vssd1 vccd1 vccd1 _09286_ sky130_fd_sc_hd__or3_1
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13855_ _06589_ _06591_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__xor2_1
XFILLER_63_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19362_ _04471_ rbzero.wall_tracer.rayAddendY\[-3\] vssd1 vssd1 vccd1 vccd1 _02851_
+ sky130_fd_sc_hd__nor2_1
X_12806_ _05539_ _05541_ _05545_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__o21ai_1
X_16574_ _09216_ vssd1 vssd1 vccd1 vccd1 _09217_ sky130_fd_sc_hd__clkbuf_4
X_10998_ _03847_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__clkbuf_1
X_13786_ _06509_ _06519_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__a21o_1
XFILLER_76_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18313_ _02011_ _02012_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__or2b_1
XFILLER_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15525_ _07981_ vssd1 vssd1 vccd1 vccd1 _08170_ sky130_fd_sc_hd__buf_4
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20178__204 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__inv_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ rbzero.debug_overlay.facingX\[-2\] rbzero.wall_tracer.rayAddendX\[6\] vssd1
+ vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__nand2_1
X_19293_ _02802_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _01827_ _01828_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__nand2_1
X_15456_ _07904_ rbzero.wall_tracer.stepDistY\[-8\] _05195_ vssd1 vssd1 vccd1 vccd1
+ _08101_ sky130_fd_sc_hd__a21o_1
XFILLER_176_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12668_ rbzero.debug_overlay.facingX\[-1\] rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__nand2_1
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14407_ _07133_ _07143_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__or2_1
XFILLER_198_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18175_ _01857_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__xnor2_1
X_11619_ rbzero.tex_r1\[47\] _04327_ _04328_ _04265_ vssd1 vssd1 vccd1 vccd1 _04398_
+ sky130_fd_sc_hd__a31o_1
X_15387_ rbzero.wall_tracer.visualWallDist\[0\] _08031_ _07904_ vssd1 vssd1 vccd1
+ vccd1 _08032_ sky130_fd_sc_hd__mux2_1
X_12599_ _05352_ _05291_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__xnor2_2
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17126_ _09757_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_144_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14338_ _07071_ _07074_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__nand2_1
XFILLER_171_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17057_ _07589_ vssd1 vssd1 vccd1 vccd1 _09697_ sky130_fd_sc_hd__inv_2
XFILLER_116_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14269_ _07005_ _06732_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__xnor2_2
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16008_ _08638_ _08651_ _08652_ vssd1 vssd1 vccd1 vccd1 _08653_ sky130_fd_sc_hd__a21oi_2
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _01454_ _01542_ _01661_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__a21oi_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20970_ clknet_leaf_3_i_clk _00739_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.vinf
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21522_ net443 _01291_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21453_ net374 _01222_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21384_ net305 _01153_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput59 net59 vssd1 vssd1 vccd1 vccd1 o_hsync sky130_fd_sc_hd__buf_2
XFILLER_153_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _04741_ _04744_ _04332_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__mux2_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10921_ _03807_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__clkbuf_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10852_ rbzero.tex_b1\[63\] net48 _03691_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__mux2_1
X_13640_ _06336_ _06375_ _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__nor3_1
XFILLER_72_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10783_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _03729_ vssd1 vssd1 vccd1 vccd1 _03735_
+ sky130_fd_sc_hd__mux2_1
X_13571_ _06306_ _06307_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__xnor2_2
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _07954_ rbzero.debug_overlay.playerY\[-4\] _05374_ vssd1 vssd1 vccd1 vccd1
+ _07955_ sky130_fd_sc_hd__mux2_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _05235_ _05276_ _05228_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or3b_1
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16290_ _08849_ _08845_ _08847_ vssd1 vssd1 vccd1 vccd1 _08935_ sky130_fd_sc_hd__and3_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15241_ rbzero.wall_tracer.wall\[0\] _03999_ _05280_ _03987_ vssd1 vssd1 vccd1 vccd1
+ _07889_ sky130_fd_sc_hd__a22o_1
XFILLER_201_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12453_ _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__buf_4
X_11404_ _04152_ _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__nor2_1
XFILLER_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12384_ net123 _05145_ _05146_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__a21oi_2
XFILLER_125_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15172_ rbzero.wall_tracer.rayAddendX\[5\] _07826_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07827_ sky130_fd_sc_hd__mux2_1
XFILLER_197_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11335_ _04101_ _04105_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__xnor2_1
X_14123_ _06851_ _06853_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__xnor2_1
XFILLER_180_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19980_ net513 _03247_ _03249_ rbzero.debug_overlay.facingY\[-2\] _03251_ vssd1 vssd1
+ vccd1 vccd1 _01022_ sky130_fd_sc_hd__a221o_1
XFILLER_207_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18931_ _02593_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__buf_4
X_11266_ gpout0.hpos\[7\] gpout0.hpos\[8\] _04045_ gpout0.hpos\[9\] vssd1 vssd1 vccd1
+ vccd1 _04046_ sky130_fd_sc_hd__a31oi_4
X_14054_ _06778_ _06790_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__xnor2_1
XFILLER_113_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13005_ _05741_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__clkbuf_4
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18862_ _02536_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__clkbuf_1
X_11197_ rbzero.map_rom.d6 _03942_ _03981_ _03985_ vssd1 vssd1 vccd1 vccd1 _03986_
+ sky130_fd_sc_hd__o31a_1
XFILLER_80_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17813_ _10130_ _10266_ _10265_ _10267_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18793_ _05204_ _02475_ _02476_ _09897_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a31o_1
XFILLER_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17744_ _01445_ _01447_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__nand2_1
X_14956_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.trackDistX\[10\] _05278_
+ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__mux2_1
XFILLER_63_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13907_ _06637_ _06619_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__and2b_1
X_17675_ _09126_ _08493_ _10238_ _10239_ vssd1 vssd1 vccd1 vccd1 _10240_ sky130_fd_sc_hd__o22ai_1
X_20062__99 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__inv_2
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14887_ _07598_ _04019_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__nand2_1
X_19414_ _02887_ _02890_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a21o_1
XFILLER_78_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16626_ _09128_ _09130_ _09131_ _09127_ vssd1 vssd1 vccd1 vccd1 _09269_ sky130_fd_sc_hd__a22o_1
X_13838_ _06258_ _06261_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__and2b_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19345_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__nand2_1
XFILLER_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16557_ _09199_ _09200_ vssd1 vssd1 vccd1 vccd1 _09201_ sky130_fd_sc_hd__xnor2_1
X_13769_ _06486_ _06487_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__or2_1
XFILLER_188_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15508_ _08131_ _08136_ _08127_ vssd1 vssd1 vccd1 vccd1 _08153_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19276_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_leak\[0\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__mux2_1
XFILLER_176_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16488_ _09127_ _09131_ vssd1 vssd1 vccd1 vccd1 _09132_ sky130_fd_sc_hd__xor2_2
X_18227_ _01925_ _01926_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__nor2_1
XFILLER_175_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15439_ _05207_ _08079_ _08082_ _08083_ vssd1 vssd1 vccd1 vccd1 _08084_ sky130_fd_sc_hd__a22o_4
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18158_ _08237_ _08493_ _08044_ _09973_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__or4_2
XFILLER_191_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17109_ _09747_ vssd1 vssd1 vccd1 vccd1 _09748_ sky130_fd_sc_hd__clkbuf_2
X_18089_ _01667_ _01676_ _01789_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__a21oi_1
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20232__253 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__inv_2
XFILLER_137_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20051_ _04990_ _04989_ _04322_ _02705_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__a41o_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20953_ clknet_leaf_95_i_clk _00722_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ clknet_leaf_88_i_clk _00653_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21505_ net426 _01274_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21436_ net357 _01205_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[15\] sky130_fd_sc_hd__dfxtp_1
X_20315__328 clknet_1_0__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__inv_2
XFILLER_148_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21367_ net288 _01136_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[10\] sky130_fd_sc_hd__dfxtp_1
X_11120_ rbzero.vga_sync.vsync vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__inv_6
XFILLER_150_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21298_ net219 _01067_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[5\] sky130_fd_sc_hd__dfxtp_1
X_11051_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _03865_ vssd1 vssd1 vccd1 vccd1 _03875_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20249_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__buf_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _05884_ _05952_ _07469_ _07538_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__a31o_1
XFILLER_92_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _08406_ _08414_ _08434_ vssd1 vssd1 vccd1 vccd1 _08435_ sky130_fd_sc_hd__a21o_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _07107_ _07350_ _07379_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__a21boi_1
XFILLER_205_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ rbzero.tex_b0\[39\] rbzero.tex_b0\[38\] _04356_ vssd1 vssd1 vccd1 vccd1 _04729_
+ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_105 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_105/HI zeros[15]
+ sky130_fd_sc_hd__conb_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_116 vssd1 vssd1 vccd1 vccd1 ones[10] top_ew_algofoogle_116/LO sky130_fd_sc_hd__conb_1
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _09906_ _10026_ vssd1 vssd1 vccd1 vccd1 _10027_ sky130_fd_sc_hd__xor2_4
X_10904_ _03798_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__clkbuf_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _07342_ _07408_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__nand2_1
X_11884_ _04241_ _04652_ _04660_ _04143_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__o211a_1
XFILLER_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16411_ _09053_ _09055_ vssd1 vssd1 vccd1 vccd1 _09056_ sky130_fd_sc_hd__xnor2_2
X_13623_ _06355_ _06359_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__xor2_1
XFILLER_60_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17391_ _09682_ _09690_ _09689_ vssd1 vssd1 vccd1 vccd1 _09958_ sky130_fd_sc_hd__a21o_2
XFILLER_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10835_ _03717_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__buf_4
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19130_ net43 rbzero.spi_registers.sclk_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02700_ sky130_fd_sc_hd__mux2_1
X_16342_ _08979_ _08986_ vssd1 vssd1 vccd1 vccd1 _08987_ sky130_fd_sc_hd__xnor2_2
XFILLER_41_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13554_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__xnor2_2
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10766_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _03718_ vssd1 vssd1 vccd1 vccd1 _03726_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19061_ rbzero.pov.spi_buffer\[61\] rbzero.pov.ready_buffer\[61\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02663_ sky130_fd_sc_hd__mux2_1
X_12505_ _05253_ _05256_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__nand3_1
X_16273_ _08816_ _08335_ _08916_ _08917_ vssd1 vssd1 vccd1 vccd1 _08918_ sky130_fd_sc_hd__o31ai_2
XFILLER_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10697_ _03689_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__clkbuf_1
X_13485_ _06211_ _06221_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18012_ _01712_ _01713_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__nor2_1
XFILLER_145_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15224_ _07873_ _07874_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__and2_1
XFILLER_185_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12436_ rbzero.wall_tracer.state\[6\] vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__buf_4
XFILLER_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15155_ rbzero.wall_tracer.rayAddendX\[4\] _07810_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07811_ sky130_fd_sc_hd__mux2_1
X_12367_ _05131_ _05132_ _05133_ _05134_ net28 _05082_ vssd1 vssd1 vccd1 vccd1 _05135_
+ sky130_fd_sc_hd__mux4_1
XFILLER_5_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14106_ _06704_ _06760_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__nor2_1
XFILLER_99_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11318_ _04060_ _04063_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__xnor2_1
X_12298_ clknet_1_1__leaf__04835_ _05046_ _05047_ vssd1 vssd1 vccd1 vccd1 _05067_
+ sky130_fd_sc_hd__and3_2
XFILLER_141_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15086_ _07741_ _07745_ _04034_ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__o21ai_1
X_19963_ rbzero.pov.ready_buffer\[37\] _03247_ _03249_ rbzero.debug_overlay.facingX\[-5\]
+ _03250_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__a221o_1
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18914_ _02580_ _02581_ _02574_ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__and3b_1
X_14037_ _06771_ _06772_ _06773_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__or3b_1
X_11249_ _04030_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__buf_2
XFILLER_141_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19894_ _07982_ _02823_ _03198_ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__o211ai_1
XFILLER_68_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18845_ _02520_ _02521_ _01908_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__a21bo_1
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18776_ _09863_ _02460_ _02461_ _09885_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__o31ai_1
X_15988_ _08008_ _08022_ vssd1 vssd1 vccd1 vccd1 _08633_ sky130_fd_sc_hd__nor2_1
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17727_ _10289_ _10291_ vssd1 vssd1 vccd1 vccd1 _10292_ sky130_fd_sc_hd__nor2_1
XFILLER_35_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14939_ _07621_ _07634_ _07635_ _07620_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__o211a_1
X_17658_ _10216_ _10221_ vssd1 vssd1 vccd1 vccd1 _10223_ sky130_fd_sc_hd__or2_1
XFILLER_91_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16609_ _08282_ _08383_ _08111_ _08570_ vssd1 vssd1 vccd1 vccd1 _09252_ sky130_fd_sc_hd__or4_1
XFILLER_63_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17589_ _10152_ _10154_ vssd1 vssd1 vccd1 vccd1 _10155_ sky130_fd_sc_hd__xor2_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19328_ net39 net38 vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__nor2_4
XFILLER_32_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19259_ _02782_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__clkbuf_4
XFILLER_177_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21221_ clknet_leaf_21_i_clk _00990_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_191_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21152_ clknet_leaf_87_i_clk _00921_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21083_ net173 _00852_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20034_ _04989_ _04037_ _02705_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__and3_1
XFILLER_86_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ clknet_leaf_93_i_clk _00705_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ clknet_leaf_5_i_clk _00636_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ _03649_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20798_ clknet_leaf_44_i_clk _00567_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10551_ _03612_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20239__259 clknet_1_0__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__inv_2
XFILLER_195_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10482_ _03576_ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__clkbuf_1
X_13270_ _05852_ _05853_ _05855_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__and3_1
XFILLER_148_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12221_ _04989_ _04990_ _04961_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__mux2_1
X_21419_ net340 _01188_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ gpout1.clk_div\[1\] _04922_ _04905_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__and3_1
XFILLER_155_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11103_ _03902_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__clkbuf_1
X_12083_ net3 net2 vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__and2_2
X_16960_ _09599_ _09600_ vssd1 vssd1 vccd1 vccd1 _09601_ sky130_fd_sc_hd__nor2_1
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15911_ _08475_ _08553_ _08554_ _08555_ vssd1 vssd1 vccd1 vccd1 _08556_ sky130_fd_sc_hd__a2bb2o_1
X_11034_ _03866_ vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__clkbuf_1
X_16891_ _08383_ _09103_ vssd1 vssd1 vccd1 vccd1 _09532_ sky130_fd_sc_hd__or2_1
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18630_ _02268_ _02284_ _02282_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a21o_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15842_ _08478_ _08485_ _08486_ vssd1 vssd1 vccd1 vccd1 _08487_ sky130_fd_sc_hd__a21o_1
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ _08445_ _09704_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__nor2_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _05208_ _08149_ vssd1 vssd1 vccd1 vccd1 _08418_ sky130_fd_sc_hd__nor2_2
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12985_ _05705_ _05708_ _05719_ _05721_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a211oi_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17512_ _10076_ _10077_ vssd1 vssd1 vccd1 vccd1 _10078_ sky130_fd_sc_hd__xor2_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _05188_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__clkbuf_4
X_18492_ _01739_ _08423_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__nor2_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ rbzero.tex_b0\[54\] _04338_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__and2_1
XFILLER_18_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17443_ _10007_ _10009_ vssd1 vssd1 vccd1 vccd1 _10010_ sky130_fd_sc_hd__xnor2_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14655_ _05742_ _05755_ _07377_ _07391_ _07375_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__a32o_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _04209_ _04639_ _04643_ _04142_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a211o_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ _06295_ _06339_ _06340_ _06342_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__a22o_1
X_17374_ _08705_ _08159_ _08151_ _09522_ vssd1 vssd1 vccd1 vccd1 _09941_ sky130_fd_sc_hd__o22a_1
X_10818_ _03753_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14586_ _07284_ _07321_ _07322_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__a21o_1
X_11798_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _04341_ vssd1 vssd1 vccd1 vccd1 _04576_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19113_ rbzero.spi_registers.mosi rbzero.spi_registers.spi_cmd\[0\] _02690_ vssd1
+ vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__mux2_1
XFILLER_201_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16325_ _08968_ _08969_ vssd1 vssd1 vccd1 vccd1 _08970_ sky130_fd_sc_hd__and2_2
X_13537_ _06225_ _06233_ _06272_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__and3_1
XFILLER_199_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10749_ _03716_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19044_ rbzero.pov.spi_buffer\[53\] rbzero.pov.ready_buffer\[53\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02654_ sky130_fd_sc_hd__mux2_1
X_16256_ _08885_ _08888_ _08900_ vssd1 vssd1 vccd1 vccd1 _08901_ sky130_fd_sc_hd__a21oi_1
XFILLER_139_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13468_ _06201_ _06204_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__xor2_1
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15207_ _07857_ _07858_ _07847_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__a21oi_1
X_12419_ net35 _05180_ _05182_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__o211a_1
X_16187_ _08829_ _08831_ vssd1 vssd1 vccd1 vccd1 _08832_ sky130_fd_sc_hd__and2b_1
X_13399_ _06132_ _06133_ _06135_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__o21ba_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15138_ _07775_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__xnor2_1
XFILLER_142_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15069_ rbzero.debug_overlay.vplaneX\[-1\] vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__clkbuf_4
X_19946_ _03236_ _03238_ _02714_ vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__o21a_1
XFILLER_114_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19877_ _02820_ _03185_ _03155_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__o21a_1
XFILLER_67_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18828_ _02503_ _02504_ _02505_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__o21a_1
X_20344__354 clknet_1_0__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__inv_2
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18759_ _02443_ _02444_ _02445_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a21oi_1
XFILLER_130_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20721_ clknet_leaf_45_i_clk _00014_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20652_ clknet_leaf_56_i_clk _00436_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20583_ rbzero.wall_tracer.rayAddendX\[-8\] _03443_ _03452_ _03453_ vssd1 vssd1 vccd1
+ vccd1 _01425_ sky130_fd_sc_hd__a22o_1
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21204_ clknet_leaf_99_i_clk _00973_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21135_ clknet_leaf_96_i_clk _00904_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21066_ net156 _00835_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_28_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20017_ _04006_ _04811_ _04813_ _03262_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__or4bb_1
XFILLER_115_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _05514_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__xnor2_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ rbzero.debug_overlay.playerY\[1\] _04449_ _04499_ rbzero.debug_overlay.playerY\[4\]
+ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__a22o_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ clknet_leaf_6_i_clk _00688_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14440_ _06680_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__and3b_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _04423_ _04426_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__and2_1
XFILLER_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10603_ rbzero.tex_g1\[53\] rbzero.tex_g1\[54\] _03635_ vssd1 vssd1 vccd1 vccd1 _03640_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14371_ _06680_ _07072_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__or2_2
XFILLER_183_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11583_ _04360_ _04361_ _04345_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__mux2_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16110_ _08741_ _08753_ _08754_ vssd1 vssd1 vccd1 vccd1 _08755_ sky130_fd_sc_hd__a21oi_1
XFILLER_122_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13322_ _05923_ _06054_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__nand2_1
XFILLER_11_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10534_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _03602_ vssd1 vssd1 vccd1 vccd1 _03604_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17090_ _09616_ _09729_ vssd1 vssd1 vccd1 vccd1 _09730_ sky130_fd_sc_hd__xnor2_2
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16041_ _08623_ _08685_ vssd1 vssd1 vccd1 vccd1 _08686_ sky130_fd_sc_hd__xnor2_1
X_10465_ _03567_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13253_ _05909_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__clkbuf_4
XFILLER_108_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12204_ _04966_ net66 _04973_ net18 vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a211o_1
XFILLER_142_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10396_ _03529_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__clkbuf_1
X_13184_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__clkinv_2
XFILLER_159_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19800_ _04867_ rbzero.pov.mosi_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1 _03129_
+ sky130_fd_sc_hd__mux2_1
X_12135_ net9 vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__inv_2
XFILLER_151_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17992_ _01687_ _01609_ _01693_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__a21oi_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03300_ clknet_0__03300_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03300_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16943_ _09445_ _09446_ vssd1 vssd1 vccd1 vccd1 _09584_ sky130_fd_sc_hd__nor2_1
X_19731_ _03093_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__clkbuf_1
X_12066_ net3 net2 vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__nor2_2
XFILLER_77_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11017_ _03857_ vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16874_ _09478_ _09479_ _09513_ vssd1 vssd1 vccd1 vccd1 _09515_ sky130_fd_sc_hd__nand3_1
X_19662_ rbzero.pov.spi_buffer\[7\] rbzero.pov.spi_buffer\[8\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03057_ sky130_fd_sc_hd__mux2_1
XFILLER_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18613_ _02307_ _02309_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__nor2_2
X_15825_ _08169_ _08469_ vssd1 vssd1 vccd1 vccd1 _08470_ sky130_fd_sc_hd__xnor2_2
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19593_ clknet_1_0__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__buf_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18544_ _02239_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__xnor2_1
X_15756_ _08108_ _08117_ vssd1 vssd1 vccd1 vccd1 _08401_ sky130_fd_sc_hd__nor2_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ _05589_ _05704_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__xnor2_2
XFILLER_79_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14707_ _07375_ _07440_ _07441_ _07443_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__a31o_1
X_18475_ _02071_ _02172_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11919_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _04271_ vssd1 vssd1 vccd1 vccd1 _04695_
+ sky130_fd_sc_hd__mux2_1
X_15687_ _05210_ _08044_ vssd1 vssd1 vccd1 vccd1 _08332_ sky130_fd_sc_hd__nor2_2
XFILLER_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12899_ _05622_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__xor2_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ _08266_ _09696_ _09989_ _09992_ vssd1 vssd1 vccd1 vccd1 _09993_ sky130_fd_sc_hd__a31oi_2
XFILLER_127_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ _05932_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__buf_2
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17357_ _09922_ _09923_ vssd1 vssd1 vccd1 vccd1 _09924_ sky130_fd_sc_hd__nand2_1
XFILLER_207_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14569_ _07305_ _07093_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__nand2_1
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16308_ _08619_ _08952_ vssd1 vssd1 vccd1 vccd1 _08953_ sky130_fd_sc_hd__xnor2_4
XFILLER_119_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17288_ _09812_ _09857_ _09858_ _09860_ vssd1 vssd1 vccd1 vccd1 _09861_ sky130_fd_sc_hd__o31ai_1
XFILLER_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19027_ rbzero.pov.spi_buffer\[45\] rbzero.pov.ready_buffer\[45\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02645_ sky130_fd_sc_hd__mux2_1
X_16239_ _08879_ _08883_ vssd1 vssd1 vccd1 vccd1 _08884_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19929_ _03223_ _03224_ _02822_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__a21oi_1
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20704_ clknet_leaf_52_i_clk _00488_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_1_0__f__03320_ clknet_0__03320_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03320_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20635_ clknet_leaf_64_i_clk _00419_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20566_ rbzero.traced_texVinit\[9\] _09764_ _07831_ _10171_ vssd1 vssd1 vccd1 vccd1
+ _01417_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20497_ rbzero.traced_texa\[2\] rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1 _03395_
+ sky130_fd_sc_hd__or2_1
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21118_ net208 _00887_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13940_ _06612_ _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__nor2_4
X_21049_ clknet_leaf_75_i_clk _00818_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13871_ _06547_ _06497_ _06498_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__and3_1
XFILLER_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15610_ _07601_ _04015_ _05198_ _08254_ vssd1 vssd1 vccd1 vccd1 _08255_ sky130_fd_sc_hd__and4_1
X_12822_ rbzero.wall_tracer.mapY\[11\] _05284_ _05533_ _05559_ vssd1 vssd1 vccd1 vccd1
+ _00418_ sky130_fd_sc_hd__a22o_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16590_ _09167_ _09174_ _09232_ vssd1 vssd1 vccd1 vccd1 _09233_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ rbzero.wall_tracer.stepDistY\[2\] vssd1 vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__inv_2
XFILLER_37_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12753_ _05204_ _05498_ _05499_ _05500_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__a31o_1
XFILLER_188_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18260_ _01952_ _01959_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__xnor2_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ rbzero.debug_overlay.facingY\[-4\] _04464_ _04465_ rbzero.debug_overlay.facingY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__a22o_1
XFILLER_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15472_ _08115_ _08116_ _08110_ vssd1 vssd1 vccd1 vccd1 _08117_ sky130_fd_sc_hd__o21a_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12684_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__or2_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ rbzero.wall_tracer.mapX\[9\] _05525_ vssd1 vssd1 vccd1 vccd1 _09793_ sky130_fd_sc_hd__nor2_1
XFILLER_129_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14423_ _07158_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__or2_1
X_18191_ _01855_ _01890_ _01891_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__nand3_1
XFILLER_202_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11635_ gpout0.hpos\[6\] _04008_ _04023_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__and3_1
XFILLER_30_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17142_ _07468_ _07544_ vssd1 vssd1 vccd1 vccd1 _09765_ sky130_fd_sc_hd__nor2_2
X_14354_ _07027_ _07029_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__nor2_1
X_11566_ _04224_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__buf_6
XFILLER_156_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20373__380 clknet_1_0__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__inv_2
XFILLER_128_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13305_ _06041_ _05940_ _05942_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__o21ai_1
X_10517_ rbzero.tex_r0\[31\] rbzero.tex_r0\[30\] _03591_ vssd1 vssd1 vccd1 vccd1 _03595_
+ sky130_fd_sc_hd__mux2_1
X_17073_ _09709_ _09712_ vssd1 vssd1 vccd1 vccd1 _09713_ sky130_fd_sc_hd__xor2_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14285_ _07020_ _07021_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__xor2_2
XFILLER_109_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11497_ rbzero.tex_r0\[14\] _04214_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__and2_1
XFILLER_170_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16024_ _08621_ _08665_ vssd1 vssd1 vccd1 vccd1 _08669_ sky130_fd_sc_hd__or2_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13236_ _05969_ _05972_ _05871_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__mux2_2
XFILLER_109_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10448_ net46 rbzero.tex_r0\[63\] _03558_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__mux2_1
XFILLER_124_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13167_ _05890_ _05903_ _05826_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__mux2_1
X_10379_ _03520_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__clkbuf_1
X_12118_ gpout0.vpos\[9\] vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__clkbuf_4
X_13098_ _05740_ _05828_ _05832_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__o211a_1
X_17975_ rbzero.wall_tracer.trackDistX\[4\] rbzero.wall_tracer.stepDistX\[4\] vssd1
+ vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__nor2_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19714_ _03084_ vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__clkbuf_1
X_16926_ _09562_ _09566_ vssd1 vssd1 vccd1 vccd1 _09567_ sky130_fd_sc_hd__xnor2_2
X_12049_ rbzero.row_render.texu\[2\] _04821_ _04822_ vssd1 vssd1 vccd1 vccd1 _04823_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03314_ _03314_ vssd1 vssd1 vccd1 vccd1 clknet_0__03314_ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19645_ _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16857_ _09487_ _09497_ vssd1 vssd1 vccd1 vccd1 _09498_ sky130_fd_sc_hd__xnor2_1
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15808_ _08452_ _08009_ vssd1 vssd1 vccd1 vccd1 _08453_ sky130_fd_sc_hd__xnor2_2
XFILLER_168_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16788_ _07579_ _07582_ vssd1 vssd1 vccd1 vccd1 _09430_ sky130_fd_sc_hd__or2_1
XFILLER_19_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15739_ _08383_ _07981_ _08180_ _08282_ vssd1 vssd1 vccd1 vccd1 _08384_ sky130_fd_sc_hd__o22ai_1
X_18527_ _02222_ _02224_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__nand2_1
XFILLER_61_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18458_ _02153_ _02154_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__and2_1
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17409_ _09288_ _09695_ vssd1 vssd1 vccd1 vccd1 _09976_ sky130_fd_sc_hd__and2_1
X_18389_ _01739_ _01475_ _01476_ _01860_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__o22ai_1
X_20420_ _03328_ _03329_ _03325_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__a21bo_1
XFILLER_146_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_7_0_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_7_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19630__82 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__inv_2
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21667_ clknet_leaf_34_i_clk _01436_ vssd1 vssd1 vccd1 vccd1 gpout4.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__03303_ clknet_0__03303_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03303_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11420_ _03475_ _04182_ _04179_ _04154_ _04199_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__a221o_1
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20618_ clknet_leaf_18_i_clk _00402_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.c6 sky130_fd_sc_hd__dfxtp_1
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21598_ net139 _01367_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ rbzero.floor_leak\[2\] _04123_ _04126_ rbzero.floor_leak\[1\] _04130_ vssd1
+ vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a221o_1
XFILLER_153_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20549_ _03430_ _03435_ _03436_ _03437_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__nand4_1
XFILLER_193_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10302_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__clkbuf_4
XFILLER_125_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14070_ _06769_ _06615_ _06738_ _06707_ _06776_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__o32ai_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] vssd1 vssd1
+ vccd1 vccd1 _04062_ sky130_fd_sc_hd__nand2_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13021_ _05710_ _05713_ _05757_ _05687_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__or4_1
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17760_ _01462_ _10205_ _01463_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__o21ba_1
X_14972_ rbzero.wall_tracer.stepDistX\[-7\] _00008_ vssd1 vssd1 vccd1 vccd1 _07656_
+ sky130_fd_sc_hd__nor2_1
XFILLER_102_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16711_ _09028_ vssd1 vssd1 vccd1 vccd1 _09353_ sky130_fd_sc_hd__inv_2
X_13923_ _06603_ _06612_ _06560_ _06601_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__o211a_1
X_17691_ _09980_ _10115_ vssd1 vssd1 vccd1 vccd1 _10256_ sky130_fd_sc_hd__or2_1
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16642_ _07575_ _08983_ _07579_ vssd1 vssd1 vccd1 vccd1 _09285_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19430_ _02912_ _02913_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__nand2_1
X_13854_ _06255_ _06265_ _06590_ vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12805_ _05539_ _05541_ _05545_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__or3_1
X_16573_ _05210_ _09215_ vssd1 vssd1 vccd1 vccd1 _09216_ sky130_fd_sc_hd__or2_1
X_19361_ rbzero.debug_overlay.vplaneY\[-7\] _02847_ vssd1 vssd1 vccd1 vccd1 _02850_
+ sky130_fd_sc_hd__nand2_1
X_13785_ _06520_ _06521_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__and2_1
X_10997_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _03843_ vssd1 vssd1 vccd1 vccd1 _03847_
+ sky130_fd_sc_hd__mux2_1
XFILLER_203_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18312_ _01915_ _01916_ _02010_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__a21o_1
X_15524_ _08120_ _08146_ _08168_ vssd1 vssd1 vccd1 vccd1 _08169_ sky130_fd_sc_hd__a21oi_2
XFILLER_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19292_ rbzero.spi_registers.new_other\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__mux2_1
X_12736_ _05461_ _05483_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__nor2_1
XFILLER_204_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _01941_ _01942_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15455_ _07933_ _07514_ _08099_ vssd1 vssd1 vccd1 vccd1 _08100_ sky130_fd_sc_hd__o21ai_2
XFILLER_203_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ _05415_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14406_ _07134_ _07135_ _07142_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__a21oi_1
X_18174_ _01858_ _01874_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__xor2_1
X_11618_ rbzero.tex_r1\[46\] _04272_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__and2_1
X_15386_ _05374_ _08030_ vssd1 vssd1 vccd1 vccd1 _08031_ sky130_fd_sc_hd__nor2_1
XFILLER_184_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12598_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__nand2_1
X_17125_ _04443_ _09750_ vssd1 vssd1 vccd1 vccd1 _09757_ sky130_fd_sc_hd__and2_1
X_14337_ _06017_ _07073_ _06770_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__a21oi_1
X_11549_ _04136_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__buf_4
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17056_ _09292_ _09695_ _08872_ vssd1 vssd1 vccd1 vccd1 _09696_ sky130_fd_sc_hd__a21oi_2
X_14268_ _07003_ _07004_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__xnor2_2
XFILLER_13_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16007_ _08639_ _08650_ vssd1 vssd1 vccd1 vccd1 _08652_ sky130_fd_sc_hd__nor2_1
X_13219_ _05740_ _05828_ _05932_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a21oi_1
XFILLER_174_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _06776_ _06610_ _06671_ _06769_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__o22a_1
XFILLER_98_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20150__179 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__inv_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17958_ _01539_ _01541_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16909_ _09539_ _09549_ vssd1 vssd1 vccd1 vccd1 _09550_ sky130_fd_sc_hd__xor2_2
XFILLER_66_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17889_ _01478_ _01480_ _01477_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a21bo_1
XFILLER_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19559_ rbzero.pov.spi_counter\[3\] _03028_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__nand2_1
XFILLER_202_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21521_ net442 _01290_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21452_ net373 _01221_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21383_ net304 _01152_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10920_ rbzero.tex_b1\[31\] rbzero.tex_b1\[32\] _03806_ vssd1 vssd1 vccd1 vccd1 _03807_
+ sky130_fd_sc_hd__mux2_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10851_ _03770_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _06107_ _06106_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__and2b_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _03734_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _05250_ _05260_ _05271_ _05275_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__o31a_1
XFILLER_200_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15240_ rbzero.wall_tracer.rayAddendX\[11\] _07855_ _07679_ _07888_ _07880_ vssd1
+ vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__a221o_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12452_ _05206_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__buf_4
XFILLER_185_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_201_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11403_ rbzero.row_render.size\[6\] _04151_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__nor2_1
XFILLER_123_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15171_ _07814_ _07815_ _04033_ _07825_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__a2bb2o_1
X_12383_ net50 _05142_ _05148_ _05149_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a211o_1
XFILLER_126_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14122_ _06822_ _06835_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__xnor2_1
X_11334_ rbzero.row_render.vinf _04113_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__nor2_8
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14053_ _06776_ _06739_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__nor2_1
X_18930_ rbzero.pov.spi_done _03480_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__nand2_1
X_11265_ _04008_ _04023_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_76_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13004_ _05740_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__buf_2
X_18861_ rbzero.wall_tracer.trackDistY\[8\] _02535_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02536_ sky130_fd_sc_hd__mux2_1
XFILLER_122_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11196_ rbzero.map_rom.f3 _03942_ _03976_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_
+ sky130_fd_sc_hd__a211o_1
X_17812_ _10110_ _09973_ _10260_ _01515_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__o31ai_2
XFILLER_95_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18792_ _02474_ _02469_ _02472_ _02473_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__a211o_1
XFILLER_121_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17743_ _01446_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
XFILLER_153_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14955_ _04019_ _07645_ _07646_ _07642_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__o211a_1
XFILLER_43_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13906_ _06640_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__inv_2
X_17674_ _08259_ vssd1 vssd1 vccd1 vccd1 _10239_ sky130_fd_sc_hd__clkbuf_4
X_14886_ rbzero.wall_tracer.visualWallDist\[-11\] vssd1 vssd1 vccd1 vccd1 _07598_
+ sky130_fd_sc_hd__inv_2
XFILLER_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19413_ _04471_ rbzero.debug_overlay.vplaneY\[-7\] vssd1 vssd1 vccd1 vccd1 _02898_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_165_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16625_ _08963_ _09119_ _09267_ vssd1 vssd1 vccd1 vccd1 _09268_ sky130_fd_sc_hd__a21bo_1
X_13837_ _06572_ _06573_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__and2_1
XFILLER_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_189_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19344_ _02828_ _02833_ _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__o21ai_1
X_16556_ _09065_ _09077_ _09078_ _09064_ vssd1 vssd1 vccd1 vccd1 _09200_ sky130_fd_sc_hd__a31o_1
X_13768_ _05825_ _06240_ _06504_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__or3_1
XFILLER_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15507_ _08135_ _08151_ vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__or2_1
X_12719_ _05430_ _05433_ _05431_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__a21boi_1
X_16487_ _09128_ _09130_ vssd1 vssd1 vccd1 vccd1 _09131_ sky130_fd_sc_hd__xor2_2
XFILLER_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19275_ _02791_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__clkbuf_4
X_13699_ _06428_ _06435_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__or2_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18226_ _01918_ _01919_ _01924_ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__and3_1
XFILLER_148_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15438_ rbzero.wall_tracer.visualWallDist\[-2\] _07925_ _05206_ vssd1 vssd1 vccd1
+ vccd1 _08083_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_129_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18157_ _01755_ _01763_ _01762_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a21bo_1
XFILLER_157_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15369_ _07913_ _07941_ _07967_ _07924_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__o22ai_1
XFILLER_11_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17108_ _03555_ _04037_ vssd1 vssd1 vccd1 vccd1 _09747_ sky130_fd_sc_hd__or2_1
X_18088_ _01667_ _01676_ _01789_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__and3_1
XFILLER_171_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17039_ _09660_ _09678_ vssd1 vssd1 vccd1 vccd1 _09679_ sky130_fd_sc_hd__xor2_2
XFILLER_132_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20050_ _03266_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__inv_2
XFILLER_113_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ clknet_leaf_2_i_clk _00721_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ clknet_leaf_88_i_clk _00652_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21504_ net425 _01273_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_158_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21435_ net356 _01204_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21366_ net287 _01135_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21297_ net218 _01066_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11050_ _03874_ vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14740_ _07107_ _07356_ _07474_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__a21oi_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11952_ _04218_ _04727_ _04253_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__o21a_1
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_106 vssd1 vssd1 vccd1 vccd1 ones[0] top_ew_algofoogle_106/LO sky130_fd_sc_hd__conb_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xtop_ew_algofoogle_117 vssd1 vssd1 vccd1 vccd1 ones[11] top_ew_algofoogle_117/LO sky130_fd_sc_hd__conb_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ rbzero.tex_b1\[39\] rbzero.tex_b1\[40\] _03795_ vssd1 vssd1 vccd1 vccd1 _03798_
+ sky130_fd_sc_hd__mux2_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _07213_ _07328_ _07332_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__a21o_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _04229_ _04655_ _04659_ _04119_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__a211o_1
XFILLER_205_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16410_ _08413_ _09054_ _08435_ vssd1 vssd1 vccd1 vccd1 _09055_ sky130_fd_sc_hd__o21a_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13622_ _06313_ _06356_ _06357_ _06358_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__o22a_1
XFILLER_60_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17390_ _09665_ _09666_ _09677_ _09956_ vssd1 vssd1 vccd1 vccd1 _09957_ sky130_fd_sc_hd__a31o_1
X_10834_ _03761_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16341_ _08239_ _08985_ vssd1 vssd1 vccd1 vccd1 _08986_ sky130_fd_sc_hd__nor2_1
X_13553_ _06112_ _06118_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__xor2_2
XFILLER_198_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10765_ _03725_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19060_ _02662_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__clkbuf_1
X_12504_ rbzero.wall_tracer.trackDistX\[0\] _05257_ _05258_ rbzero.wall_tracer.trackDistX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__o22a_1
X_16272_ _08215_ _08226_ _08135_ _08160_ vssd1 vssd1 vccd1 vccd1 _08917_ sky130_fd_sc_hd__or4_1
XFILLER_73_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ _06219_ _06220_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__and2_1
XFILLER_186_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10696_ rbzero.tex_g1\[9\] rbzero.tex_g1\[10\] _03680_ vssd1 vssd1 vccd1 vccd1 _03689_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18011_ _01710_ _01711_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__and2_1
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15223_ _07872_ _07868_ _07869_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__or3_1
XFILLER_200_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12435_ _05194_ _03914_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__nor2_1
XFILLER_172_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15154_ _04034_ _07799_ _07807_ _07809_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__a22o_1
X_12366_ _04891_ _04992_ _04890_ _04892_ _05091_ _05083_ vssd1 vssd1 vccd1 vccd1 _05134_
+ sky130_fd_sc_hd__mux4_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14105_ _06703_ _06841_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__xnor2_2
X_11317_ _04075_ _04093_ _04096_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__o21a_1
XFILLER_180_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15085_ _07743_ _07744_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__nor2_1
X_19962_ _02695_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__buf_6
XFILLER_99_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12297_ _05062_ _05064_ _05065_ _05047_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a2bb2o_1
X_18913_ rbzero.spi_registers.spi_counter\[1\] rbzero.spi_registers.spi_counter\[0\]
+ _02558_ rbzero.spi_registers.spi_counter\[2\] vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a31o_1
X_14036_ _06009_ _06658_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__nor2_1
X_11248_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__buf_2
XFILLER_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19893_ rbzero.pov.ready_buffer\[45\] _02823_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__nand2_1
XFILLER_110_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18844_ _02517_ _02518_ _02519_ _09807_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__o31a_1
XFILLER_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11179_ _03957_ _03965_ _03966_ _03967_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__and4b_2
XFILLER_110_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18775_ _02457_ _02458_ _02459_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15987_ _08630_ _08631_ vssd1 vssd1 vccd1 vccd1 _08632_ sky130_fd_sc_hd__xor2_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17726_ _10039_ _10163_ _10290_ vssd1 vssd1 vccd1 vccd1 _10291_ sky130_fd_sc_hd__a21oi_1
XFILLER_76_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14938_ rbzero.wall_tracer.visualWallDist\[4\] _07618_ vssd1 vssd1 vccd1 vccd1 _07635_
+ sky130_fd_sc_hd__or2_1
XFILLER_169_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17657_ _10216_ _10221_ vssd1 vssd1 vccd1 vccd1 _10222_ sky130_fd_sc_hd__and2_1
XFILLER_24_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14869_ _07394_ _07440_ _07441_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__and3_1
XFILLER_51_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ _09248_ _09250_ vssd1 vssd1 vccd1 vccd1 _09251_ sky130_fd_sc_hd__and2_1
XFILLER_35_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17588_ _09972_ _10010_ _10153_ vssd1 vssd1 vccd1 vccd1 _10154_ sky130_fd_sc_hd__a21boi_1
XFILLER_204_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19327_ rbzero.spi_registers.got_new_vshift _02730_ _02728_ _02813_ vssd1 vssd1 vccd1
+ vccd1 _00803_ sky130_fd_sc_hd__a31o_1
X_16539_ _09156_ _09182_ vssd1 vssd1 vccd1 vccd1 _09183_ sky130_fd_sc_hd__xnor2_2
XFILLER_52_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19258_ _02772_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__or3b_1
XFILLER_104_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18209_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.stepDistX\[6\] vssd1
+ vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__and2_1
X_19189_ rbzero.floor_leak\[5\] _02732_ _02739_ _02722_ vssd1 vssd1 vccd1 vccd1 _00745_
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21220_ clknet_leaf_20_i_clk _00989_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[-9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_172_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20156__185 clknet_1_1__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__inv_2
XFILLER_132_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21151_ clknet_leaf_87_i_clk _00920_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21082_ net172 _00851_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20033_ _09753_ _03267_ _03274_ _03272_ _04884_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__a32o_1
XFILLER_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ clknet_leaf_92_i_clk _00704_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20321__333 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__inv_2
XFILLER_54_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20866_ clknet_leaf_94_i_clk _00635_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20797_ clknet_leaf_43_i_clk _00566_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ rbzero.tex_r0\[15\] rbzero.tex_r0\[14\] _03602_ vssd1 vssd1 vccd1 vccd1 _03612_
+ sky130_fd_sc_hd__mux2_1
XFILLER_195_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10481_ rbzero.tex_r0\[48\] rbzero.tex_r0\[47\] _03569_ vssd1 vssd1 vccd1 vccd1 _03576_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12220_ gpout0.vpos\[5\] vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__buf_2
XFILLER_136_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21418_ net339 _01187_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ _04906_ _04909_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nor2_1
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21349_ net270 _01118_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11102_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _03898_ vssd1 vssd1 vccd1 vccd1 _03902_
+ sky130_fd_sc_hd__mux2_1
XFILLER_190_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12082_ net51 _04837_ net47 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a21o_1
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15910_ _08008_ _07967_ vssd1 vssd1 vccd1 vccd1 _08555_ sky130_fd_sc_hd__nor2_1
XFILLER_2_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11033_ rbzero.tex_b0\[42\] rbzero.tex_b0\[41\] _03865_ vssd1 vssd1 vccd1 vccd1 _03866_
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16890_ _09529_ _09530_ vssd1 vssd1 vccd1 vccd1 _09531_ sky130_fd_sc_hd__xnor2_2
XFILLER_76_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _08137_ _08143_ vssd1 vssd1 vccd1 vccd1 _08486_ sky130_fd_sc_hd__xnor2_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ _02167_ _02255_ _02256_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a21o_1
XFILLER_58_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _05208_ _08157_ vssd1 vssd1 vccd1 vccd1 _08417_ sky130_fd_sc_hd__nor2_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _05596_ _05720_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__xor2_4
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17511_ _09526_ _08427_ vssd1 vssd1 vccd1 vccd1 _10077_ sky130_fd_sc_hd__nor2_1
XFILLER_166_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11935_ _04709_ _04710_ _04247_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__mux2_1
X_14723_ _07456_ _07458_ _07459_ vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__mux2_1
X_18491_ _02187_ _02188_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__nand2_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _09692_ _09717_ _10008_ vssd1 vssd1 vccd1 vccd1 _10009_ sky130_fd_sc_hd__a21o_2
X_14654_ _05741_ _07383_ _07390_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__a21oi_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11866_ _04640_ _04641_ _04642_ _04139_ _04253_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__o221a_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20296__310 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__inv_2
XFILLER_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13605_ _06292_ _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__xnor2_1
X_10817_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _03751_ vssd1 vssd1 vccd1 vccd1 _03753_
+ sky130_fd_sc_hd__mux2_1
X_17373_ _09664_ _09665_ vssd1 vssd1 vccd1 vccd1 _09940_ sky130_fd_sc_hd__nand2_1
X_14585_ _07279_ _07282_ _07281_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__o21bai_1
X_11797_ _04573_ _04574_ _04217_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__mux2_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19112_ rbzero.spi_registers.spi_counter\[3\] rbzero.spi_registers.spi_counter\[2\]
+ _02567_ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__or4_2
X_16324_ _08959_ _08967_ vssd1 vssd1 vccd1 vccd1 _08969_ sky130_fd_sc_hd__or2_1
X_13536_ _06225_ _06233_ _06272_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10748_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _03706_ vssd1 vssd1 vccd1 vccd1 _03716_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16255_ _08892_ _08899_ vssd1 vssd1 vccd1 vccd1 _08900_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19043_ _02653_ vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13467_ _06160_ _06202_ _06203_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__a21o_1
XFILLER_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10679_ _03646_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__clkbuf_4
X_15206_ _07821_ _07742_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__or2_1
X_12418_ net37 _05184_ _05145_ net34 vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__and4bb_1
XFILLER_127_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16186_ _08788_ _08830_ vssd1 vssd1 vccd1 vccd1 _08831_ sky130_fd_sc_hd__nand2_1
XFILLER_138_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13398_ _06065_ _06058_ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__nor3_1
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15137_ _07791_ _07793_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__xnor2_1
X_12349_ net29 net28 _05116_ net30 vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a31o_1
XFILLER_142_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15068_ rbzero.debug_overlay.vplaneX\[-1\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__or2_1
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19945_ rbzero.pov.ready_buffer\[58\] _03164_ _03197_ _03237_ vssd1 vssd1 vccd1 vccd1
+ _03238_ sky130_fd_sc_hd__o211a_1
XFILLER_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14019_ _06752_ _06754_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__and2_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19876_ rbzero.debug_overlay.playerX\[4\] _03180_ vssd1 vssd1 vccd1 vccd1 _03185_
+ sky130_fd_sc_hd__and2b_1
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18827_ _02503_ _02504_ _02505_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__nor3_1
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18758_ _02443_ _02444_ _02445_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__and3_1
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17709_ _10123_ _10148_ _10145_ vssd1 vssd1 vccd1 vccd1 _10274_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18689_ _02252_ _02286_ _02384_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a21oi_1
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20720_ clknet_leaf_59_i_clk _00010_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20651_ clknet_leaf_56_i_clk _00435_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20582_ _07688_ _07831_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__nor2_1
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21203_ clknet_leaf_98_i_clk _00972_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21134_ clknet_leaf_96_i_clk _00903_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21065_ net155 _00834_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20016_ _03474_ _04809_ _03554_ _04815_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__nor4_1
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _04022_ _04444_ _04440_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__and3_1
X_20918_ clknet_leaf_6_i_clk _00687_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _04008_ _04023_ _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a21oi_4
XFILLER_199_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20849_ clknet_leaf_45_i_clk _00618_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10602_ _03639_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14370_ _05893_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__clkbuf_4
XFILLER_168_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11582_ rbzero.tex_r1\[23\] rbzero.tex_r1\[22\] _04290_ vssd1 vssd1 vccd1 vccd1 _04361_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13321_ _06053_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a21o_1
X_10533_ _03603_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16040_ _07923_ _08125_ vssd1 vssd1 vccd1 vccd1 _08685_ sky130_fd_sc_hd__nor2_1
X_13252_ _05939_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__clkinv_2
X_10464_ rbzero.tex_r0\[56\] rbzero.tex_r0\[55\] _03558_ vssd1 vssd1 vccd1 vccd1 _03567_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12203_ _04966_ _04325_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__nor2_1
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13183_ _05834_ _05913_ _05914_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__a31o_2
X_10395_ rbzero.tex_r1\[22\] rbzero.tex_r1\[23\] _03527_ vssd1 vssd1 vccd1 vccd1 _03529_
+ sky130_fd_sc_hd__mux2_1
XFILLER_163_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12134_ net11 net10 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__nor2_2
X_17991_ _01691_ _01692_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__nand2_1
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19730_ rbzero.pov.spi_buffer\[39\] rbzero.pov.spi_buffer\[40\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03093_ sky130_fd_sc_hd__mux2_1
X_12065_ net7 net6 vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__nor2_2
X_16942_ _09517_ _09582_ vssd1 vssd1 vccd1 vccd1 _09583_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11016_ rbzero.tex_b0\[50\] rbzero.tex_b0\[49\] _03854_ vssd1 vssd1 vccd1 vccd1 _03857_
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20328__339 clknet_1_0__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__inv_2
X_19661_ _03056_ vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16873_ _09478_ _09479_ _09513_ vssd1 vssd1 vccd1 vccd1 _09514_ sky130_fd_sc_hd__a21o_1
XFILLER_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18612_ _02218_ _02220_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__o21a_1
XFILLER_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ _08439_ _08468_ vssd1 vssd1 vccd1 vccd1 _08469_ sky130_fd_sc_hd__xor2_2
XFILLER_93_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ _01620_ _09292_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__nor2_1
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15755_ _08372_ _08399_ vssd1 vssd1 vccd1 vccd1 _08400_ sky130_fd_sc_hd__xor2_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12967_ _05591_ _05593_ _05628_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__o21a_1
XFILLER_206_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _07375_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__nor2_1
X_11918_ _04345_ _04693_ _04253_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__o21a_1
X_18474_ _08257_ _09027_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__nor2_1
X_15686_ _08039_ vssd1 vssd1 vccd1 vccd1 _08331_ sky130_fd_sc_hd__buf_4
X_12898_ _05609_ _05619_ _05562_ _05566_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__o211a_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _08873_ _09977_ _09991_ _08872_ vssd1 vssd1 vccd1 vccd1 _09992_ sky130_fd_sc_hd__o22a_1
XFILLER_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11849_ _04620_ _04622_ _04625_ _04306_ _04241_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__a221o_1
XFILLER_33_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14637_ _05741_ _07348_ _07353_ _07373_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__a31o_1
XFILLER_127_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17356_ _08335_ _09483_ _09910_ vssd1 vssd1 vccd1 vccd1 _09923_ sky130_fd_sc_hd__o21ai_1
X_14568_ _07297_ _07299_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__xor2_1
XFILLER_202_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16307_ _08950_ _08946_ _08671_ vssd1 vssd1 vccd1 vccd1 _08952_ sky130_fd_sc_hd__a21o_1
X_13519_ _05921_ _06176_ _06215_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__and3_1
X_14499_ _07188_ _07189_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__xor2_1
X_17287_ _09807_ _09859_ vssd1 vssd1 vccd1 vccd1 _09860_ sky130_fd_sc_hd__or2_1
XFILLER_118_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19026_ _02644_ vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__clkbuf_1
X_20073__109 clknet_1_0__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__inv_2
X_16238_ _08881_ _08882_ vssd1 vssd1 vccd1 vccd1 _08883_ sky130_fd_sc_hd__xor2_1
XFILLER_133_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16169_ _08791_ _08787_ _08790_ vssd1 vssd1 vccd1 vccd1 _08814_ sky130_fd_sc_hd__a21oi_1
XFILLER_142_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19928_ rbzero.debug_overlay.playerY\[1\] _03216_ rbzero.debug_overlay.playerY\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__o21ai_1
XFILLER_69_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19859_ rbzero.debug_overlay.playerX\[1\] _03167_ vssd1 vssd1 vccd1 vccd1 _03171_
+ sky130_fd_sc_hd__nor2_1
XFILLER_68_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20268__286 clknet_1_1__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__inv_2
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_3_0_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20703_ clknet_leaf_52_i_clk _00487_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_93_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20634_ clknet_leaf_12_i_clk _00418_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20565_ rbzero.traced_texVinit\[8\] _09764_ _07831_ _10027_ vssd1 vssd1 vccd1 vccd1
+ _01416_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_165_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20496_ _09750_ _03392_ _03394_ _03250_ rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1
+ _01397_ sky130_fd_sc_hd__a32o_1
XFILLER_124_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21117_ net207 _00886_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21048_ clknet_leaf_75_i_clk _00817_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13870_ _06552_ _06606_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__and2_2
X_12821_ _05557_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12752_ _03926_ _05394_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__nor2_1
X_15540_ _07894_ _05456_ _08184_ _05193_ vssd1 vssd1 vccd1 vccd1 _08185_ sky130_fd_sc_hd__a211o_2
XFILLER_15_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11703_ rbzero.debug_overlay.facingY\[-6\] _04475_ _04458_ rbzero.debug_overlay.facingY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a22o_1
X_15471_ _08097_ _08042_ vssd1 vssd1 vccd1 vccd1 _08116_ sky130_fd_sc_hd__or2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ rbzero.debug_overlay.facingX\[-5\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__nand2_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _07114_ _07127_ _07157_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__a21oi_1
X_17210_ rbzero.wall_tracer.mapX\[9\] _05525_ vssd1 vssd1 vccd1 vccd1 _09792_ sky130_fd_sc_hd__and2_1
X_11634_ _04206_ _04412_ _04314_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a21o_1
X_18190_ _01887_ _01888_ _01889_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__a21o_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17141_ rbzero.row_render.size\[4\] _09762_ _07541_ _07756_ vssd1 vssd1 vccd1 vccd1
+ _00532_ sky130_fd_sc_hd__a22o_1
X_14353_ _07044_ _07089_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__xnor2_1
X_11565_ rbzero.tex_r1\[7\] rbzero.tex_r1\[6\] _04342_ vssd1 vssd1 vccd1 vccd1 _04344_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13304_ _05846_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__buf_2
X_10516_ _03594_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__clkbuf_1
X_17072_ _09710_ _09566_ _09711_ vssd1 vssd1 vccd1 vccd1 _09712_ sky130_fd_sc_hd__a21oi_4
XFILLER_155_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14284_ _06766_ _06767_ _06782_ _06781_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__a31o_1
X_11496_ _04274_ _04275_ _04226_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__mux2_1
XFILLER_143_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13235_ _05800_ _05864_ _05970_ _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__o211a_1
X_16023_ _08658_ _08662_ _08667_ vssd1 vssd1 vccd1 vccd1 _08668_ sky130_fd_sc_hd__o21a_2
XFILLER_115_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10447_ _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13166_ _05783_ _05757_ _05791_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__mux2_1
X_10378_ rbzero.tex_r1\[30\] rbzero.tex_r1\[31\] _03516_ vssd1 vssd1 vccd1 vccd1 _03520_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12117_ gpout0.vpos\[4\] gpout0.vpos\[5\] _04840_ vssd1 vssd1 vccd1 vccd1 _04889_
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17974_ _05203_ _01674_ _01676_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__or3b_2
X_13097_ _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__clkbuf_4
X_19616__69 clknet_1_0__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__inv_2
X_19713_ net512 rbzero.pov.spi_buffer\[32\] _03081_ vssd1 vssd1 vccd1 vccd1 _03084_
+ sky130_fd_sc_hd__mux2_1
X_16925_ _08816_ _09565_ vssd1 vssd1 vccd1 vccd1 _09566_ sky130_fd_sc_hd__nor2_2
X_12048_ rbzero.row_render.texu\[3\] _03473_ _04163_ vssd1 vssd1 vccd1 vccd1 _04822_
+ sky130_fd_sc_hd__or3b_1
XFILLER_78_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03313_ _03313_ vssd1 vssd1 vccd1 vccd1 clknet_0__03313_ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19644_ _03046_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__buf_4
X_16856_ _09495_ _09496_ vssd1 vssd1 vccd1 vccd1 _09497_ sky130_fd_sc_hd__nor2_1
XFILLER_20_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15807_ _08010_ _07997_ vssd1 vssd1 vccd1 vccd1 _08452_ sky130_fd_sc_hd__nand2_1
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16787_ _08230_ rbzero.wall_tracer.stepDistY\[9\] vssd1 vssd1 vccd1 vccd1 _09429_
+ sky130_fd_sc_hd__nand2_1
X_13999_ _06719_ _06723_ _06734_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__and3_1
XFILLER_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18526_ _02223_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__inv_2
XFILLER_179_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15738_ _08276_ vssd1 vssd1 vccd1 vccd1 _08383_ sky130_fd_sc_hd__clkbuf_4
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18457_ _02153_ _02154_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__nor2_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15669_ _07913_ _07996_ _07932_ _07924_ vssd1 vssd1 vccd1 vccd1 _08314_ sky130_fd_sc_hd__o22ai_1
X_17408_ _09553_ _09974_ _09687_ _09684_ vssd1 vssd1 vccd1 vccd1 _09975_ sky130_fd_sc_hd__a22o_1
X_18388_ _01739_ _01860_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__or4_1
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17339_ _09594_ _09596_ _09737_ _09905_ vssd1 vssd1 vccd1 vccd1 _09906_ sky130_fd_sc_hd__a31oi_4
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20274__290 clknet_1_1__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__inv_2
XFILLER_162_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19009_ _02635_ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21666_ clknet_leaf_34_i_clk _01435_ vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__03302_ clknet_0__03302_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03302_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20617_ clknet_leaf_8_i_clk _00401_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.d6 sky130_fd_sc_hd__dfxtp_2
X_21597_ net138 _01366_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11350_ rbzero.floor_leak\[1\] _04125_ _04129_ rbzero.floor_leak\[0\] vssd1 vssd1
+ vccd1 vccd1 _04130_ sky130_fd_sc_hd__o211a_1
X_20548_ _03435_ _03436_ _03437_ _03430_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__a22o_1
XFILLER_119_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10301_ gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__inv_2
XFILLER_153_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11281_ rbzero.traced_texVinit\[6\] rbzero.spi_registers.vshift\[3\] vssd1 vssd1
+ vccd1 vccd1 _04061_ sky130_fd_sc_hd__or2_1
X_20479_ _03373_ _03377_ _03378_ _03379_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__o211a_1
XFILLER_180_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13020_ _05584_ _05714_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__xnor2_2
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14971_ _00008_ _07514_ _07655_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16710_ _08162_ _09351_ vssd1 vssd1 vccd1 vccd1 _09352_ sky130_fd_sc_hd__or2_1
XFILLER_120_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13922_ _05825_ _06658_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__nor2_2
XFILLER_48_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17690_ _08767_ _09693_ vssd1 vssd1 vccd1 vccd1 _10255_ sky130_fd_sc_hd__nor2_1
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ _09283_ rbzero.wall_tracer.stepDistY\[8\] vssd1 vssd1 vccd1 vccd1 _09284_
+ sky130_fd_sc_hd__nand2_1
XFILLER_63_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13853_ _06219_ _06266_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__nor2_1
XFILLER_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19360_ rbzero.debug_overlay.vplaneY\[-7\] _02847_ vssd1 vssd1 vccd1 vccd1 _02849_
+ sky130_fd_sc_hd__or2_1
X_12804_ rbzero.wall_tracer.mapY\[8\] _05404_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__xor2_1
X_16572_ rbzero.wall_tracer.visualWallDist\[8\] _04015_ vssd1 vssd1 vccd1 vccd1 _09215_
+ sky130_fd_sc_hd__nand2_4
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10996_ _03846_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__clkbuf_1
X_13784_ _06509_ _06519_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__xor2_1
X_18311_ _01915_ _01916_ _02010_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__and3_1
XFILLER_203_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15523_ _08154_ _08167_ vssd1 vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__xor2_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19291_ _02800_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__buf_4
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12735_ _05466_ _05468_ _05469_ _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__or4_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20104__138 clknet_1_1__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__inv_2
XFILLER_31_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _08275_ _09217_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__or2_1
XFILLER_176_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _07971_ _05481_ _08098_ vssd1 vssd1 vccd1 vccd1 _08099_ sky130_fd_sc_hd__o21ai_2
X_12666_ rbzero.map_rom.f4 _05410_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__mux2_1
XFILLER_187_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11617_ rbzero.tex_r1\[45\] rbzero.tex_r1\[44\] _04392_ vssd1 vssd1 vccd1 vccd1 _04396_
+ sky130_fd_sc_hd__mux2_1
X_14405_ _07140_ _07141_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__and2b_1
XFILLER_198_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18173_ _01865_ _01873_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12597_ _05350_ _05293_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__xor2_1
X_15385_ rbzero.debug_overlay.playerY\[-1\] rbzero.debug_overlay.playerY\[-2\] _08029_
+ vssd1 vssd1 vccd1 vccd1 _08030_ sky130_fd_sc_hd__or3_1
XFILLER_11_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17124_ _04422_ _09748_ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__nor2_1
XFILLER_129_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11548_ _04135_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__buf_4
X_14336_ _06776_ _07072_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__or2_1
XFILLER_128_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17055_ _05210_ rbzero.wall_tracer.stepDistX\[8\] vssd1 vssd1 vccd1 vccd1 _09695_
+ sky130_fd_sc_hd__nand2_4
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14267_ _06744_ _06751_ _06755_ vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__a21oi_2
XFILLER_7_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11479_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _04213_ vssd1 vssd1 vccd1 vccd1 _04259_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13218_ _05952_ _05916_ _05954_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16006_ _08639_ _08650_ vssd1 vssd1 vccd1 vccd1 _08651_ sky130_fd_sc_hd__xor2_1
X_14198_ _06769_ _06610_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__nor2_1
XFILLER_87_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _05884_ _05885_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__nor2_1
XFILLER_97_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _01572_ _01659_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16908_ _09547_ _09548_ vssd1 vssd1 vccd1 vccd1 _09549_ sky130_fd_sc_hd__and2b_1
X_17888_ _01580_ _01590_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__xor2_1
XFILLER_39_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16839_ _09351_ vssd1 vssd1 vccd1 vccd1 _09480_ sky130_fd_sc_hd__clkbuf_4
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19558_ _03028_ _03029_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__nor2_1
X_18509_ _02067_ _02069_ _02066_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__o21ba_1
XFILLER_94_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19489_ _02948_ _02954_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__nand2_1
XFILLER_90_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21520_ net441 _01289_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20079__115 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__inv_2
XFILLER_194_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21451_ net372 _01220_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21382_ net303 _01151_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10850_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _03762_ vssd1 vssd1 vccd1 vccd1 _03770_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ rbzero.tex_g0\[34\] rbzero.tex_g0\[33\] _03729_ vssd1 vssd1 vccd1 vccd1 _03734_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ rbzero.wall_tracer.trackDistY\[3\] _05264_ _05269_ _05274_ vssd1 vssd1 vccd1
+ vccd1 _05275_ sky130_fd_sc_hd__a22o_1
XFILLER_200_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _05195_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__buf_4
XFILLER_184_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21649_ clknet_leaf_41_i_clk _01418_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_20290__305 clknet_1_1__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__inv_2
XFILLER_184_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11402_ rbzero.row_render.size\[7\] _04152_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15170_ _07823_ _07824_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__and2b_1
XFILLER_197_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12382_ net34 vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__inv_2
XFILLER_123_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14121_ _06699_ _06855_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__xnor2_1
X_11333_ _04110_ _04112_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__xnor2_2
XFILLER_10_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14052_ _06787_ _06788_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11264_ gpout0.vpos\[9\] gpout0.vpos\[8\] gpout0.vpos\[7\] net1 vssd1 vssd1 vccd1
+ vccd1 _04044_ sky130_fd_sc_hd__or4b_1
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13003_ _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__clkbuf_2
XFILLER_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18860_ _02128_ _02130_ _02533_ _02534_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a22o_1
X_11195_ _03919_ _03925_ rbzero.map_rom.a6 _03983_ rbzero.map_rom.f1 vssd1 vssd1 vccd1
+ vccd1 _03984_ sky130_fd_sc_hd__a2111o_1
XFILLER_122_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17811_ _10115_ _01514_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__nand2_1
XFILLER_121_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ _02472_ _02473_ _02474_ _02469_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__o211ai_1
X_17742_ _08331_ _09610_ _10201_ _10200_ _09368_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__o32a_1
X_14954_ rbzero.wall_tracer.visualWallDist\[9\] _07594_ vssd1 vssd1 vccd1 vccd1 _07646_
+ sky130_fd_sc_hd__or2_1
XFILLER_47_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ _06595_ _06598_ _06640_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__a21o_2
X_17673_ _08044_ vssd1 vssd1 vccd1 vccd1 _10238_ sky130_fd_sc_hd__clkbuf_4
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14885_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.trackDistX\[-11\]
+ _07592_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__mux2_1
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19412_ _02893_ _02894_ _02895_ _02879_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a22o_1
X_16624_ _08383_ _09114_ _09121_ vssd1 vssd1 vccd1 vccd1 _09267_ sky130_fd_sc_hd__or3_1
X_13836_ _06242_ _06244_ _06571_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__nand3_1
XFILLER_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19343_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__nand2_1
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16555_ _09197_ _09198_ vssd1 vssd1 vccd1 vccd1 _09199_ sky130_fd_sc_hd__or2b_1
X_10979_ _03837_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__clkbuf_1
X_13767_ _06501_ _06503_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__and2_1
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15506_ _08150_ vssd1 vssd1 vccd1 vccd1 _08151_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12718_ _05463_ _05465_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__xnor2_2
X_19274_ rbzero.spi_registers.spi_cmd\[0\] _02772_ rbzero.spi_registers.spi_cmd\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__or3b_1
X_16486_ _08242_ _09129_ _08170_ vssd1 vssd1 vccd1 vccd1 _09130_ sky130_fd_sc_hd__a21oi_2
XFILLER_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13698_ _06431_ _06433_ _06434_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__o21a_1
XFILLER_148_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18225_ _01918_ _01919_ _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15437_ _07951_ _08081_ vssd1 vssd1 vccd1 vccd1 _08082_ sky130_fd_sc_hd__nand2_1
X_12649_ _05388_ _05399_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__nand2_1
XFILLER_175_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18156_ _01743_ _01750_ _01856_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__a21o_1
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15368_ _08011_ _07969_ vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__xor2_1
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17107_ rbzero.wall_tracer.texu\[5\] _09085_ _04035_ _09746_ vssd1 vssd1 vccd1 vccd1
+ _00516_ sky130_fd_sc_hd__o211a_1
XFILLER_156_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14319_ _07007_ _07012_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__nand2_1
X_18087_ _01788_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__inv_2
X_15299_ _07942_ _07943_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__nand2_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17038_ _09667_ _09677_ vssd1 vssd1 vccd1 vccd1 _09678_ sky130_fd_sc_hd__xor2_2
XFILLER_144_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ rbzero.pov.spi_buffer\[27\] rbzero.pov.ready_buffer\[27\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02625_ sky130_fd_sc_hd__mux2_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20951_ clknet_leaf_2_i_clk _00720_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20882_ clknet_leaf_98_i_clk _00651_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21503_ net424 _01272_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21434_ net355 _01203_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21365_ net286 _01134_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20316_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__buf_1
XFILLER_163_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21296_ net217 _01065_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20133__164 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__inv_2
XFILLER_153_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ rbzero.tex_b0\[35\] rbzero.tex_b0\[34\] _04262_ vssd1 vssd1 vccd1 vccd1 _04727_
+ sky130_fd_sc_hd__mux2_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xtop_ew_algofoogle_107 vssd1 vssd1 vccd1 vccd1 ones[1] top_ew_algofoogle_107/LO sky130_fd_sc_hd__conb_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _03797_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__clkbuf_1
Xtop_ew_algofoogle_118 vssd1 vssd1 vccd1 vccd1 ones[12] top_ew_algofoogle_118/LO sky130_fd_sc_hd__conb_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11882_ _04139_ _04656_ _04657_ _04658_ _04208_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__o221a_1
X_14670_ _07218_ _07323_ _07345_ _07334_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__and4_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13621_ _05920_ _06009_ _06310_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__o21a_1
X_10833_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _03751_ vssd1 vssd1 vccd1 vccd1 _03761_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16340_ _08980_ _08984_ _08147_ vssd1 vssd1 vccd1 vccd1 _08985_ sky130_fd_sc_hd__a21o_1
X_10764_ rbzero.tex_g0\[42\] rbzero.tex_g0\[41\] _03718_ vssd1 vssd1 vccd1 vccd1 _03725_
+ sky130_fd_sc_hd__mux2_1
X_13552_ _06286_ _06288_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__or2_1
XFILLER_9_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ rbzero.wall_tracer.trackDistY\[-1\] vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__inv_2
XFILLER_201_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16271_ _08215_ _08162_ _08160_ _08226_ vssd1 vssd1 vccd1 vccd1 _08916_ sky130_fd_sc_hd__o22a_1
X_13483_ _06212_ _06213_ _06218_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__or3_1
XFILLER_200_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10695_ _03688_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__clkbuf_1
X_18010_ _01710_ _01711_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__nor2_1
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15222_ _07868_ _07869_ _07872_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__o21ai_1
X_12434_ _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__buf_4
XFILLER_173_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12365_ _04989_ _04990_ _05083_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__mux2_1
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15153_ _04033_ _07808_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__nor2_1
XFILLER_154_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14104_ _06818_ _06840_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__xor2_2
X_11316_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__inv_2
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15084_ _07742_ rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _07744_
+ sky130_fd_sc_hd__and2_1
X_19961_ _03248_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__clkbuf_4
X_12296_ net45 _05043_ _05049_ gpout3.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _05065_
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18912_ rbzero.spi_registers.spi_counter\[2\] rbzero.spi_registers.spi_counter\[1\]
+ rbzero.spi_registers.spi_counter\[0\] _02558_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__and4_1
X_14035_ _05984_ _06769_ _06658_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__a21o_1
XFILLER_180_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11247_ _04003_ _03913_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__nor2_1
XFILLER_171_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19892_ _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__buf_2
XFILLER_79_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18843_ _02517_ _02518_ _02519_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__o21ai_1
X_11178_ rbzero.othery\[1\] _03942_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__xnor2_1
XFILLER_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18774_ _02457_ _02458_ _02459_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__and3_1
XFILLER_110_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15986_ _07988_ _07964_ _07965_ vssd1 vssd1 vccd1 vccd1 _08631_ sky130_fd_sc_hd__or3_1
XFILLER_83_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17725_ _10160_ _10162_ vssd1 vssd1 vccd1 vccd1 _10290_ sky130_fd_sc_hd__nor2_1
X_14937_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.trackDistX\[4\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__mux2_1
XFILLER_36_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17656_ _10219_ _10220_ vssd1 vssd1 vccd1 vccd1 _10221_ sky130_fd_sc_hd__and2_1
X_14868_ _07583_ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16607_ _09249_ _08356_ _09247_ vssd1 vssd1 vccd1 vccd1 _09250_ sky130_fd_sc_hd__o21ai_1
X_13819_ _06333_ _06377_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__nor2_1
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17587_ _10007_ _10009_ vssd1 vssd1 vccd1 vccd1 _10153_ sky130_fd_sc_hd__or2b_1
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14799_ _07487_ _07456_ _07529_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__a21oi_4
X_19326_ _02819_ vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__clkbuf_1
X_16538_ _09158_ _09181_ vssd1 vssd1 vccd1 vccd1 _09182_ sky130_fd_sc_hd__xnor2_2
XFILLER_17_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19257_ rbzero.spi_registers.got_new_sky _02730_ _02728_ _02781_ vssd1 vssd1 vccd1
+ vccd1 _00771_ sky130_fd_sc_hd__a31o_1
X_16469_ _09090_ _09112_ vssd1 vssd1 vccd1 vccd1 _09113_ sky130_fd_sc_hd__xor2_2
XFILLER_192_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18208_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.stepDistX\[6\] vssd1
+ vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__nor2_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19188_ rbzero.spi_registers.new_leak\[5\] _02733_ vssd1 vssd1 vccd1 vccd1 _02739_
+ sky130_fd_sc_hd__or2_1
XFILLER_191_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18139_ _01740_ _01742_ _01738_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a21bo_1
XFILLER_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21150_ clknet_leaf_86_i_clk _00919_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21081_ net171 _00850_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20032_ _02705_ _03273_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__nor2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_60_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20934_ clknet_leaf_78_i_clk _00703_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19585__41 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__inv_2
XFILLER_54_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20865_ clknet_leaf_95_i_clk _00634_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_75_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20796_ clknet_leaf_42_i_clk _00565_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10480_ _03575_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21417_ net338 _01186_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12150_ net11 net10 _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__and3b_1
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21348_ net269 _01117_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11101_ _03901_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_i_clk clknet_opt_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12081_ net3 _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__and2_1
X_21279_ clknet_leaf_95_i_clk _01048_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_done
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11032_ _03717_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__clkbuf_4
XFILLER_77_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _08479_ _08484_ vssd1 vssd1 vccd1 vccd1 _08485_ sky130_fd_sc_hd__or2b_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _08124_ vssd1 vssd1 vccd1 vccd1 _08416_ sky130_fd_sc_hd__inv_2
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12983_ _05563_ _05566_ _05594_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__and3_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _10073_ _10075_ vssd1 vssd1 vccd1 vccd1 _10076_ sky130_fd_sc_hd__nand2_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14722_ _05871_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__buf_4
X_18490_ _01860_ _01475_ _01476_ _09141_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__o22ai_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _04263_ vssd1 vssd1 vccd1 vccd1 _04710_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _09714_ _09716_ vssd1 vssd1 vccd1 vccd1 _10008_ sky130_fd_sc_hd__nor2_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ _05741_ _07389_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__nor2_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ rbzero.tex_g1\[1\] rbzero.tex_g1\[0\] _04336_ vssd1 vssd1 vccd1 vccd1 _04642_
+ sky130_fd_sc_hd__mux2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _05877_ _05923_ _06116_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__and3_1
X_17372_ _09641_ _09644_ _09643_ vssd1 vssd1 vccd1 vccd1 _09939_ sky130_fd_sc_hd__a21bo_1
X_10816_ _03752_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__clkbuf_1
X_11796_ rbzero.tex_g0\[41\] rbzero.tex_g0\[40\] _04341_ vssd1 vssd1 vccd1 vccd1 _04574_
+ sky130_fd_sc_hd__mux2_1
X_14584_ _07304_ _07308_ _07315_ _07318_ _07320_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__a41o_1
XFILLER_198_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19111_ _02557_ _02558_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__nand2_1
XFILLER_203_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16323_ _08959_ _08967_ vssd1 vssd1 vccd1 vccd1 _08968_ sky130_fd_sc_hd__nand2_1
XFILLER_186_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13535_ _06269_ _06271_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__xor2_1
X_10747_ _03715_ vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19042_ rbzero.pov.spi_buffer\[52\] rbzero.pov.ready_buffer\[52\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02653_ sky130_fd_sc_hd__mux2_1
X_16254_ _08897_ _08898_ vssd1 vssd1 vccd1 vccd1 _08899_ sky130_fd_sc_hd__nor2_1
X_10678_ _03679_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__clkbuf_1
X_13466_ _05974_ _06159_ _06161_ _05983_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__o22a_1
X_15205_ _07821_ _07742_ vssd1 vssd1 vccd1 vccd1 _07857_ sky130_fd_sc_hd__nand2_1
X_12417_ _05146_ _04738_ _05183_ net35 net36 vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__o2111a_1
XFILLER_173_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16185_ _07981_ _08128_ vssd1 vssd1 vccd1 vccd1 _08830_ sky130_fd_sc_hd__nor2_1
X_13397_ _06084_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__clkbuf_4
XFILLER_86_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15136_ _07777_ _07792_ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__or2_1
XFILLER_5_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12348_ _03473_ _04814_ _04317_ _04809_ _05083_ _05082_ vssd1 vssd1 vccd1 vccd1 _05116_
+ sky130_fd_sc_hd__mux4_1
XFILLER_154_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12279_ net42 _05046_ _05047_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__and3_1
X_15067_ _07679_ vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__buf_4
X_19944_ _03235_ _03920_ _03227_ _02822_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__a31o_1
XFILLER_142_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ _06752_ _06754_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nor2_1
XFILLER_68_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19875_ _03138_ _03183_ rbzero.debug_overlay.playerX\[4\] vssd1 vssd1 vccd1 vccd1
+ _03184_ sky130_fd_sc_hd__o21a_1
X_18826_ _02498_ _02500_ _02497_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__a21boi_1
XFILLER_83_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18757_ _02435_ _02437_ _02436_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__o21bai_1
X_15969_ _08585_ _08613_ vssd1 vssd1 vccd1 vccd1 _08614_ sky130_fd_sc_hd__nand2_1
XFILLER_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17708_ _10264_ _10272_ vssd1 vssd1 vccd1 vccd1 _10273_ sky130_fd_sc_hd__xnor2_2
X_18688_ _02254_ _02285_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__and2_1
XFILLER_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17639_ _10202_ _10203_ vssd1 vssd1 vccd1 vccd1 _10204_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20650_ clknet_leaf_56_i_clk _00434_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19309_ _02810_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20581_ _07687_ _07686_ _07685_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__a21bo_1
XFILLER_143_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21202_ clknet_leaf_98_i_clk _00971_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.sclk_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21133_ clknet_leaf_95_i_clk _00902_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21064_ net154 _00833_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20015_ _03257_ _03258_ _03261_ _03209_ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__o211a_1
XFILLER_115_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20245__265 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__inv_2
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20917_ clknet_leaf_6_i_clk _00686_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ _04005_ _04023_ gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__a21oi_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ clknet_leaf_48_i_clk _00617_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ rbzero.tex_g1\[54\] rbzero.tex_g1\[55\] _03635_ vssd1 vssd1 vccd1 vccd1 _03639_
+ sky130_fd_sc_hd__mux2_1
X_11581_ rbzero.tex_r1\[21\] rbzero.tex_r1\[20\] _04290_ vssd1 vssd1 vccd1 vccd1 _04360_
+ sky130_fd_sc_hd__mux2_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20779_ clknet_leaf_72_i_clk _00548_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10532_ rbzero.tex_r0\[24\] rbzero.tex_r0\[23\] _03602_ vssd1 vssd1 vccd1 vccd1 _03603_
+ sky130_fd_sc_hd__mux2_1
X_13320_ _05947_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__clkbuf_4
XFILLER_156_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10463_ _03566_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__clkbuf_1
X_13251_ _05941_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__clkbuf_4
XFILLER_202_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12202_ net19 vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__inv_2
XFILLER_182_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13182_ _05814_ _05915_ _05918_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a21oi_1
XFILLER_164_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10394_ _03528_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12133_ net12 net13 vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__nor2_2
XFILLER_159_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ _01688_ _01690_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__or2_1
X_12064_ net5 net4 vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__or2_1
X_16941_ _09579_ _09581_ vssd1 vssd1 vccd1 vccd1 _09582_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11015_ _03856_ vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19660_ rbzero.pov.spi_buffer\[6\] rbzero.pov.spi_buffer\[7\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03056_ sky130_fd_sc_hd__mux2_1
X_16872_ _09498_ _09512_ vssd1 vssd1 vccd1 vccd1 _09513_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18611_ _02215_ _02217_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__or2_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ _08464_ _08466_ _08467_ vssd1 vssd1 vccd1 vccd1 _08468_ sky130_fd_sc_hd__a21oi_2
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18542_ _02237_ _02238_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__xnor2_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _08391_ _08397_ _08398_ vssd1 vssd1 vccd1 vccd1 _08399_ sky130_fd_sc_hd__a21oi_2
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12966_ _05701_ _05702_ _05683_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__nor3_4
XFILLER_79_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _05894_ _07041_ _07389_ _05741_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__a22o_1
X_18473_ _02169_ _02170_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__xnor2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11917_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _04290_ vssd1 vssd1 vccd1 vccd1 _04693_
+ sky130_fd_sc_hd__mux2_1
X_15685_ _08035_ _08046_ _08329_ _08104_ vssd1 vssd1 vccd1 vccd1 _08330_ sky130_fd_sc_hd__or4_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _05626_ _05633_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__xor2_2
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17424_ _09990_ vssd1 vssd1 vccd1 vccd1 _09991_ sky130_fd_sc_hd__clkbuf_4
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14636_ _05779_ _07362_ _07372_ _05892_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__o211a_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _04623_ _04624_ _04304_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__mux2_1
XFILLER_199_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _08335_ _09483_ _09910_ vssd1 vssd1 vccd1 vccd1 _09922_ sky130_fd_sc_hd__or3_1
X_14567_ _07302_ _07303_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__nor2_1
XFILLER_186_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11779_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _04262_ vssd1 vssd1 vccd1 vccd1 _04557_
+ sky130_fd_sc_hd__mux2_1
XFILLER_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16306_ _08944_ _08948_ _08949_ _08950_ vssd1 vssd1 vccd1 vccd1 _08951_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_119_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13518_ _06154_ _06205_ _06254_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__a21bo_1
XFILLER_186_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17286_ _09061_ _09062_ vssd1 vssd1 vccd1 vccd1 _09859_ sky130_fd_sc_hd__nand2_2
XFILLER_201_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14498_ _07227_ _07231_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__xor2_1
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19025_ rbzero.pov.spi_buffer\[44\] rbzero.pov.ready_buffer\[44\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02644_ sky130_fd_sc_hd__mux2_1
X_16237_ _08857_ _08859_ _08855_ vssd1 vssd1 vccd1 vccd1 _08882_ sky130_fd_sc_hd__a21boi_1
X_13449_ _06175_ _06185_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16168_ _08791_ _08787_ _08790_ vssd1 vssd1 vccd1 vccd1 _08813_ sky130_fd_sc_hd__and3_1
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15119_ _04462_ rbzero.debug_overlay.vplaneX\[-7\] _07774_ _07775_ vssd1 vssd1 vccd1
+ vccd1 _07777_ sky130_fd_sc_hd__nor4_1
XFILLER_141_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16099_ _08704_ _08706_ vssd1 vssd1 vccd1 vccd1 _08744_ sky130_fd_sc_hd__xnor2_2
XFILLER_173_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19927_ rbzero.debug_overlay.playerY\[2\] rbzero.debug_overlay.playerY\[1\] _03216_
+ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__or3_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19858_ rbzero.debug_overlay.playerX\[0\] _03139_ _03170_ net60 vssd1 vssd1 vccd1
+ vccd1 _00983_ sky130_fd_sc_hd__a211o_1
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18809_ rbzero.wall_tracer.trackDistY\[1\] _02490_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02491_ sky130_fd_sc_hd__mux2_1
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19642__92 clknet_1_1__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__inv_2
X_19789_ _03123_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03289_ clknet_0__03289_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03289_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20702_ clknet_leaf_52_i_clk _00486_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20633_ clknet_leaf_13_i_clk _00417_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20564_ rbzero.traced_texVinit\[7\] _03443_ _09771_ _09739_ vssd1 vssd1 vccd1 vccd1
+ _01415_ sky130_fd_sc_hd__a22o_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20495_ _03393_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__inv_2
XFILLER_121_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21116_ net206 _00885_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21047_ clknet_leaf_76_i_clk _00816_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20169__196 clknet_1_1__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__inv_2
XFILLER_47_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12820_ rbzero.wall_tracer.mapY\[11\] _05404_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ rbzero.map_rom.f4 _05497_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__nand2_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _04040_ _04315_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__or2_1
X_15470_ _08110_ _08114_ vssd1 vssd1 vccd1 vccd1 _08115_ sky130_fd_sc_hd__nand2_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _05422_ _05423_ _05428_ _05429_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__o31ai_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _07114_ _07127_ _07157_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__and3_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ rbzero.color_sky\[1\] rbzero.color_floor\[1\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04412_ sky130_fd_sc_hd__mux2_1
XFILLER_196_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _07536_ _09763_ rbzero.row_render.size\[3\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00531_ sky130_fd_sc_hd__a2bb2o_1
X_14352_ _07086_ _07088_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__xor2_1
X_11564_ rbzero.tex_r1\[5\] rbzero.tex_r1\[4\] _04342_ vssd1 vssd1 vccd1 vccd1 _04343_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ _06033_ _06036_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__nand2_1
X_10515_ rbzero.tex_r0\[32\] rbzero.tex_r0\[31\] _03591_ vssd1 vssd1 vccd1 vccd1 _03594_
+ sky130_fd_sc_hd__mux2_1
X_17071_ _09560_ _09561_ vssd1 vssd1 vccd1 vccd1 _09711_ sky130_fd_sc_hd__nor2_1
X_11495_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _04273_ vssd1 vssd1 vccd1 vccd1 _04275_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14283_ _07017_ _07019_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__xor2_2
XFILLER_171_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16022_ _08657_ _08656_ vssd1 vssd1 vccd1 vccd1 _08667_ sky130_fd_sc_hd__or2b_1
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10446_ _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__buf_4
X_13234_ _05725_ _05764_ _05793_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__mux2_1
XFILLER_196_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10377_ _03519_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__clkbuf_1
X_13165_ _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__inv_2
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12116_ _04886_ _04887_ _04840_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__mux2_1
X_17973_ _01669_ _01675_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__or2_1
X_13096_ _05700_ _05703_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__or2_1
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12047_ _04814_ _03473_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__nand2_1
X_16924_ _09283_ rbzero.wall_tracer.stepDistY\[10\] _08235_ _09564_ vssd1 vssd1 vccd1
+ vccd1 _09565_ sky130_fd_sc_hd__a22oi_4
X_19712_ _03083_ vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03312_ _03312_ vssd1 vssd1 vccd1 vccd1 clknet_0__03312_ sky130_fd_sc_hd__clkbuf_16
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16855_ _09492_ _09494_ vssd1 vssd1 vccd1 vccd1 _09496_ sky130_fd_sc_hd__and2_1
X_19643_ _03020_ _03019_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__nand2_1
XFILLER_38_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15806_ _08444_ _08450_ vssd1 vssd1 vccd1 vccd1 _08451_ sky130_fd_sc_hd__xor2_2
X_16786_ _09426_ _09427_ vssd1 vssd1 vccd1 vccd1 _09428_ sky130_fd_sc_hd__xnor2_2
XFILLER_207_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13998_ _06719_ _06723_ _06734_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__a21oi_2
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18525_ _02138_ _02120_ _02221_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__and3_2
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15737_ _08375_ _08381_ vssd1 vssd1 vccd1 vccd1 _08382_ sky130_fd_sc_hd__xor2_1
XFILLER_34_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12949_ _05582_ _05600_ _05628_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__o21a_1
XFILLER_207_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18456_ _10248_ _09991_ _02046_ _02045_ _10266_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__o32a_1
XFILLER_34_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15668_ _08298_ _08312_ vssd1 vssd1 vccd1 vccd1 _08313_ sky130_fd_sc_hd__xor2_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17407_ _08895_ _09973_ vssd1 vssd1 vccd1 vccd1 _09974_ sky130_fd_sc_hd__nor2_1
XFILLER_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14619_ _07354_ _07355_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__nor2_1
X_18387_ _02085_ _01985_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__nand2_1
X_15599_ _08183_ _08185_ _07602_ _08230_ _05208_ vssd1 vssd1 vccd1 vccd1 _08244_ sky130_fd_sc_hd__a2111o_1
XFILLER_18_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17338_ _09592_ _09904_ _09736_ vssd1 vssd1 vccd1 vccd1 _09905_ sky130_fd_sc_hd__a21o_1
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17269_ _09812_ _09841_ _09842_ _09843_ vssd1 vssd1 vccd1 vccd1 _09844_ sky130_fd_sc_hd__o31ai_1
XFILLER_134_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19008_ rbzero.pov.spi_buffer\[36\] rbzero.pov.ready_buffer\[36\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02635_ sky130_fd_sc_hd__mux2_1
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20386__12 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__inv_2
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03301_ clknet_0__03301_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03301_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21665_ clknet_leaf_34_i_clk _01434_ vssd1 vssd1 vccd1 vccd1 gpout3.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20357__366 clknet_1_1__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__inv_2
XFILLER_138_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20616_ clknet_leaf_71_i_clk _00012_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[2\]
+ sky130_fd_sc_hd__dfxtp_4
X_21596_ net137 _01365_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20547_ rbzero.traced_texa\[9\] rbzero.texV\[9\] _03432_ vssd1 vssd1 vccd1 vccd1
+ _03437_ sky130_fd_sc_hd__a21o_1
XFILLER_138_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10300_ gpout0.hpos\[7\] vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__buf_4
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ rbzero.texV\[7\] _04059_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__xor2_1
X_20478_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 _03379_
+ sky130_fd_sc_hd__nand2_1
XFILLER_192_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14970_ rbzero.wall_tracer.stepDistX\[-8\] _00008_ vssd1 vssd1 vccd1 vccd1 _07655_
+ sky130_fd_sc_hd__nor2_1
XFILLER_102_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13921_ _06615_ _06641_ _06642_ _06657_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__a31o_4
XFILLER_75_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16640_ _08230_ vssd1 vssd1 vccd1 vccd1 _09283_ sky130_fd_sc_hd__buf_6
X_13852_ _06568_ _06588_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12803_ _05533_ _05542_ _05544_ _05284_ rbzero.wall_tracer.mapY\[7\] vssd1 vssd1
+ vccd1 vccd1 _00414_ sky130_fd_sc_hd__a32o_1
XFILLER_90_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16571_ _09212_ _09213_ vssd1 vssd1 vccd1 vccd1 _09214_ sky130_fd_sc_hd__nand2_1
X_13783_ _06432_ _06504_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__xnor2_1
XFILLER_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10995_ rbzero.tex_b0\[60\] rbzero.tex_b0\[59\] _03843_ vssd1 vssd1 vccd1 vccd1 _03846_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18310_ _01917_ _02009_ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__xor2_1
XFILLER_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15522_ _08165_ _08166_ vssd1 vssd1 vccd1 vccd1 _08167_ sky130_fd_sc_hd__nor2_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19290_ rbzero.spi_registers.spi_done _03480_ _02569_ vssd1 vssd1 vccd1 vccd1 _02800_
+ sky130_fd_sc_hd__and3_1
X_12734_ _05472_ _05475_ _05478_ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__or4_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18241_ _01939_ _01940_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__xnor2_2
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _07893_ _05353_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _08098_
+ sky130_fd_sc_hd__o21a_1
X_12665_ _05413_ vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__buf_6
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14404_ _07122_ _07124_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__xnor2_1
X_18172_ _01870_ _01872_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__xor2_1
X_11616_ _04393_ _04394_ _04304_ vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__mux2_1
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15384_ rbzero.debug_overlay.playerY\[-3\] _07952_ vssd1 vssd1 vccd1 vccd1 _08029_
+ sky130_fd_sc_hd__or2_1
X_12596_ _05294_ _05290_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__and2b_1
XFILLER_184_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17123_ _09756_ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14335_ _06658_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__buf_2
X_11547_ rbzero.tex_r1\[14\] _04213_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__and2_1
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17054_ _08873_ _09693_ vssd1 vssd1 vccd1 vccd1 _09694_ sky130_fd_sc_hd__nor2_2
X_14266_ _07001_ _07002_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__or2_2
XFILLER_109_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11478_ _04226_ _04257_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__or2_1
XFILLER_48_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16005_ _08640_ _08648_ _08649_ vssd1 vssd1 vccd1 vccd1 _08650_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13217_ _05952_ _05953_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__nor2_1
X_10429_ _03546_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14197_ _06929_ _06933_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__nand2_1
XFILLER_125_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _05713_ _05718_ _05721_ _05715_ _05778_ _05801_ vssd1 vssd1 vccd1 vccd1 _05885_
+ sky130_fd_sc_hd__mux4_1
XFILLER_174_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17956_ _01656_ _01658_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _05642_ _05636_ _05791_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__mux2_1
XFILLER_85_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16907_ _09418_ _09422_ _09546_ _09542_ vssd1 vssd1 vccd1 vccd1 _09548_ sky130_fd_sc_hd__a211o_1
X_17887_ _01588_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__nor2_1
X_19626_ clknet_1_1__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__buf_1
X_16838_ _09404_ _09383_ vssd1 vssd1 vccd1 vccd1 _09479_ sky130_fd_sc_hd__or2b_1
XFILLER_20_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16769_ _09270_ _09409_ _09410_ vssd1 vssd1 vccd1 vccd1 _09411_ sky130_fd_sc_hd__a21o_1
X_19557_ rbzero.pov.spi_counter\[2\] _03022_ _03020_ vssd1 vssd1 vccd1 vccd1 _03029_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_20_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18508_ _02100_ _02062_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__or2b_1
XFILLER_34_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19488_ _02904_ rbzero.wall_tracer.rayAddendY\[6\] vssd1 vssd1 vccd1 vccd1 _02968_
+ sky130_fd_sc_hd__xor2_1
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18439_ _02131_ _02137_ rbzero.wall_tracer.trackDistX\[8\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00597_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21450_ net371 _01219_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21381_ net302 _01150_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20194_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__buf_1
XFILLER_27_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _03733_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12450_ rbzero.debug_overlay.playerY\[0\] _03925_ _05204_ vssd1 vssd1 vccd1 vccd1
+ _05205_ sky130_fd_sc_hd__mux2_1
XFILLER_200_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21648_ clknet_leaf_45_i_clk _01417_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11401_ rbzero.row_render.size\[9\] _04153_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__and2_1
XFILLER_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12381_ net52 _05144_ _05139_ net49 _05147_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a221o_1
X_21579_ net500 _01348_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_80 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14120_ _06820_ _06838_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11332_ _04049_ _04111_ vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14051_ _06777_ _06778_ _06779_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__a21bo_1
X_11263_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] _04042_ vssd1 vssd1 vccd1
+ vccd1 _04043_ sky130_fd_sc_hd__or4_1
XFILLER_107_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13002_ _05700_ _05732_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__or3b_1
X_11194_ rbzero.map_rom.f4 rbzero.map_rom.d6 _03982_ _03924_ vssd1 vssd1 vccd1 vccd1
+ _03983_ sky130_fd_sc_hd__a22o_1
XFILLER_161_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17810_ _09292_ _09695_ _08767_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__a21oi_2
XFILLER_122_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18790_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__nand2_1
XFILLER_122_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20110__143 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__inv_2
X_17741_ _10204_ _10213_ _10211_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a21o_1
X_14953_ rbzero.wall_tracer.trackDistY\[9\] rbzero.wall_tracer.trackDistX\[9\] _05278_
+ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__mux2_1
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13904_ _06595_ _06598_ _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__nand3_4
X_17672_ _08259_ _09126_ _08493_ _08044_ vssd1 vssd1 vccd1 vccd1 _10237_ sky130_fd_sc_hd__or4_1
XFILLER_48_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14884_ _07591_ _07593_ _07596_ _04039_ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__o211a_1
XFILLER_90_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16623_ _09240_ _09265_ vssd1 vssd1 vccd1 vccd1 _09266_ sky130_fd_sc_hd__xnor2_1
X_19411_ _02879_ _02893_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__nand4_2
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13835_ _06242_ _06244_ _06571_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__a21o_1
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19342_ _02829_ _02832_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__and2_1
X_16554_ _09194_ _09196_ vssd1 vssd1 vccd1 vccd1 _09198_ sky130_fd_sc_hd__nand2_1
X_13766_ _05855_ _06153_ _06501_ _06502_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__nand4_1
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10978_ rbzero.tex_b1\[3\] rbzero.tex_b1\[4\] _03828_ vssd1 vssd1 vccd1 vccd1 _03837_
+ sky130_fd_sc_hd__mux2_1
XFILLER_206_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15505_ _08147_ _08149_ vssd1 vssd1 vccd1 vccd1 _08150_ sky130_fd_sc_hd__or2_2
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ _05421_ _05430_ _05433_ _05464_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__a31o_1
X_19273_ rbzero.spi_registers.got_new_floor _02730_ _02728_ _02790_ vssd1 vssd1 vccd1
+ vccd1 _00778_ sky130_fd_sc_hd__a31o_1
X_16485_ _05209_ rbzero.wall_tracer.stepDistX\[4\] vssd1 vssd1 vccd1 vccd1 _09129_
+ sky130_fd_sc_hd__nand2_2
XFILLER_203_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13697_ _06429_ _06430_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__or2b_1
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18224_ _01922_ _01923_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__nand2_1
XFILLER_15_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15436_ _08080_ rbzero.debug_overlay.playerY\[-2\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _08081_ sky130_fd_sc_hd__mux2_2
XFILLER_50_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12648_ _05389_ _05392_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__or2_1
XFILLER_129_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18155_ _01748_ _01749_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__nor2_1
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15367_ _07969_ _08011_ vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__or2b_1
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12579_ _05320_ _05322_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__and3_1
XFILLER_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17106_ _05194_ _09744_ _09745_ vssd1 vssd1 vccd1 vccd1 _09746_ sky130_fd_sc_hd__or3b_1
XFILLER_8_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14318_ _07053_ _07054_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__or2_1
XFILLER_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18086_ _01786_ _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__nor2_1
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15298_ _07913_ _07932_ _07941_ _07924_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__o22ai_1
XFILLER_102_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17037_ _09673_ _09676_ vssd1 vssd1 vccd1 vccd1 _09677_ sky130_fd_sc_hd__xor2_2
XFILLER_132_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14249_ _06909_ _06985_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__nand2_1
XFILLER_172_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _02624_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__clkbuf_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _01639_ _01640_ _01635_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a21o_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20085__120 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__inv_2
X_20950_ clknet_leaf_2_i_clk _00719_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_96_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20881_ clknet_leaf_97_i_clk _00650_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21502_ net423 _01271_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21433_ net354 _01202_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21364_ net285 _01133_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21295_ net216 _01064_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_104_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _04345_ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__or2_1
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ rbzero.tex_b1\[40\] rbzero.tex_b1\[41\] _03795_ vssd1 vssd1 vccd1 vccd1 _03797_
+ sky130_fd_sc_hd__mux2_1
Xtop_ew_algofoogle_108 vssd1 vssd1 vccd1 vccd1 ones[2] top_ew_algofoogle_108/LO sky130_fd_sc_hd__conb_1
XFILLER_205_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_119 vssd1 vssd1 vccd1 vccd1 ones[13] top_ew_algofoogle_119/LO sky130_fd_sc_hd__conb_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ rbzero.tex_g1\[30\] _04342_ _04126_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__a21o_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13620_ _05990_ _06016_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__or2_1
XFILLER_199_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10832_ _03760_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13551_ _05988_ _06287_ _06286_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__nor3_1
XFILLER_41_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10763_ _03724_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12502_ rbzero.wall_tracer.trackDistY\[0\] vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__inv_2
X_16270_ _08863_ _08914_ vssd1 vssd1 vccd1 vccd1 _08915_ sky130_fd_sc_hd__or2_1
XFILLER_40_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13482_ _06212_ _06213_ _06218_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__o21ai_2
XFILLER_41_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ rbzero.tex_g1\[10\] rbzero.tex_g1\[11\] _03680_ vssd1 vssd1 vccd1 vccd1 _03688_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15221_ _07870_ _07871_ vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__and2_1
X_12433_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__clkinv_4
XFILLER_166_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15152_ _07804_ _07806_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__and2_1
X_12364_ _04886_ _04887_ _05083_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__mux2_1
XFILLER_148_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ _06820_ _06838_ _06839_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__a21oi_2
X_11315_ _04069_ _04094_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__or2_1
XFILLER_154_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15083_ _07742_ rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _07743_
+ sky130_fd_sc_hd__nor2_1
X_19960_ _02708_ _03137_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__nand2_4
X_12295_ net50 _05043_ _05063_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18911_ _02579_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__clkbuf_1
X_14034_ _06002_ _06770_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__and2_1
X_11246_ _04029_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__clkbuf_4
XFILLER_122_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19891_ net39 _03137_ _02708_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__o21a_1
XFILLER_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18842_ _02510_ _02512_ _02511_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__a21boi_1
XFILLER_122_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11177_ rbzero.othery\[0\] rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18773_ _02450_ _02453_ _02451_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__o21ai_1
X_15985_ _07980_ _07938_ _07939_ vssd1 vssd1 vccd1 vccd1 _08630_ sky130_fd_sc_hd__or3_1
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17724_ _10186_ _10288_ vssd1 vssd1 vccd1 vccd1 _10289_ sky130_fd_sc_hd__xnor2_1
X_14936_ _07621_ _07632_ _07633_ _07620_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__o211a_1
XFILLER_76_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17655_ _09522_ _08427_ _10218_ vssd1 vssd1 vccd1 vccd1 _10220_ sky130_fd_sc_hd__o21ai_1
XFILLER_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14867_ rbzero.wall_tracer.stepDistY\[9\] _07582_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07583_ sky130_fd_sc_hd__mux2_1
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16606_ _09243_ vssd1 vssd1 vccd1 vccd1 _09249_ sky130_fd_sc_hd__clkbuf_4
X_13818_ _06464_ _06552_ _06554_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__a21bo_1
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17586_ _10109_ _10151_ vssd1 vssd1 vccd1 vccd1 _10152_ sky130_fd_sc_hd__xnor2_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14798_ _07486_ _07433_ _07442_ _07528_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__a31o_1
XFILLER_189_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16537_ _09160_ _09180_ vssd1 vssd1 vccd1 vccd1 _09181_ sky130_fd_sc_hd__xnor2_1
X_19325_ rbzero.spi_registers.new_vshift\[5\] rbzero.spi_registers.spi_buffer\[5\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__mux2_1
X_13749_ _06483_ _06485_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__xor2_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16468_ _09110_ _09111_ vssd1 vssd1 vccd1 vccd1 _09112_ sky130_fd_sc_hd__nor2_1
X_19256_ _02774_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__inv_2
XFILLER_176_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18207_ _01906_ _01907_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__or2_1
X_15419_ _08056_ _08063_ vssd1 vssd1 vccd1 vccd1 _08064_ sky130_fd_sc_hd__xor2_1
X_19187_ rbzero.floor_leak\[4\] _02732_ _02738_ _02722_ vssd1 vssd1 vccd1 vccd1 _00744_
+ sky130_fd_sc_hd__o211a_1
XFILLER_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16399_ _09030_ _09043_ vssd1 vssd1 vccd1 vccd1 _09044_ sky130_fd_sc_hd__xnor2_1
XFILLER_163_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18138_ _01719_ _01721_ _01718_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__a21bo_1
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18069_ _01768_ _01769_ _01753_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a21o_1
X_20117__149 clknet_1_0__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__inv_2
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21080_ net170 _00849_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_171_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20031_ _04884_ _02704_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__nor2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20933_ clknet_leaf_78_i_clk _00702_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20864_ clknet_leaf_95_i_clk _00633_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20795_ clknet_leaf_46_i_clk _00564_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21416_ net337 _01185_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21347_ net268 _01116_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11100_ rbzero.tex_b0\[10\] rbzero.tex_b0\[9\] _03898_ vssd1 vssd1 vccd1 vccd1 _03901_
+ sky130_fd_sc_hd__mux2_1
XFILLER_190_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12080_ net2 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__clkinv_2
XFILLER_151_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21278_ clknet_leaf_78_i_clk _01047_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_89_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11031_ _03864_ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15770_ _08059_ _08334_ _08335_ vssd1 vssd1 vccd1 vccd1 _08415_ sky130_fd_sc_hd__or3_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12982_ _05716_ _05718_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__or2_1
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14721_ _07403_ _07457_ _07433_ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__mux2_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ rbzero.tex_b0\[49\] rbzero.tex_b0\[48\] _04263_ vssd1 vssd1 vccd1 vccd1 _04709_
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _09986_ _10006_ vssd1 vssd1 vccd1 vccd1 _10007_ sky130_fd_sc_hd__xnor2_2
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ _07386_ _07388_ _05931_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__mux2_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ rbzero.tex_g1\[2\] _04356_ _04126_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__a21o_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20222__244 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__inv_2
X_13603_ _06065_ _05940_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__nor2_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17371_ _09936_ _09937_ vssd1 vssd1 vccd1 vccd1 _09938_ sky130_fd_sc_hd__and2_1
X_10815_ rbzero.tex_g0\[18\] rbzero.tex_g0\[17\] _03751_ vssd1 vssd1 vccd1 vccd1 _03752_
+ sky130_fd_sc_hd__mux2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14583_ _07316_ _07319_ _07317_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__a21oi_1
X_11795_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _04211_ vssd1 vssd1 vccd1 vccd1 _04573_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16322_ _08961_ _08966_ vssd1 vssd1 vccd1 vccd1 _08967_ sky130_fd_sc_hd__xor2_1
X_19110_ _02688_ vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__clkbuf_1
X_13534_ _06211_ _06221_ _06270_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__a21oi_1
X_10746_ rbzero.tex_g0\[50\] rbzero.tex_g0\[49\] _03706_ vssd1 vssd1 vccd1 vccd1 _03715_
+ sky130_fd_sc_hd__mux2_1
XFILLER_203_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19041_ _02652_ vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__clkbuf_1
X_16253_ _08896_ _08893_ _08894_ vssd1 vssd1 vccd1 vccd1 _08898_ sky130_fd_sc_hd__and3_1
XFILLER_9_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13465_ _05974_ _06161_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__nor2_1
XFILLER_201_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10677_ rbzero.tex_g1\[18\] rbzero.tex_g1\[19\] _03669_ vssd1 vssd1 vccd1 vccd1 _03679_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15204_ _07756_ _07845_ _07846_ _07856_ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__a31o_1
X_12416_ _05146_ net64 vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__nand2_1
XFILLER_185_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16184_ _08170_ _08042_ _08128_ _08180_ vssd1 vssd1 vccd1 vccd1 _08829_ sky130_fd_sc_hd__o22a_1
XFILLER_12_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13396_ _06065_ _06080_ _06084_ _06057_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__o22a_1
XFILLER_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15135_ _07778_ _07779_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__nor2_1
X_12347_ _05090_ _05102_ _05110_ _05114_ net30 vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__a221oi_2
XFILLER_153_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15066_ _07727_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__clkbuf_1
X_19943_ _03235_ _03233_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__nor2_1
X_12278_ net23 net22 vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__nor2_1
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14017_ _06753_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__inv_2
X_11229_ _04013_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__buf_4
X_19874_ _02820_ _03180_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__nor2_1
XFILLER_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18825_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] vssd1
+ vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__and2_1
XFILLER_68_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18756_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.stepDistY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__nand2_1
XFILLER_110_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15968_ _08609_ _08611_ _08612_ vssd1 vssd1 vccd1 vccd1 _08613_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17707_ _10126_ _10269_ _10271_ vssd1 vssd1 vccd1 vccd1 _10272_ sky130_fd_sc_hd__a21oi_2
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14919_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.trackDistX\[-2\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__mux2_1
X_18687_ _02305_ _02306_ _02303_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__o21ba_1
X_15899_ _08511_ _08543_ vssd1 vssd1 vccd1 vccd1 _08544_ sky130_fd_sc_hd__xor2_4
XFILLER_24_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17638_ _08037_ _09704_ vssd1 vssd1 vccd1 vccd1 _10203_ sky130_fd_sc_hd__nor2_1
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17569_ _10134_ _10130_ _10131_ _10132_ vssd1 vssd1 vccd1 vccd1 _10135_ sky130_fd_sc_hd__a31o_1
X_20197__221 clknet_1_0__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__inv_2
XFILLER_17_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19308_ rbzero.spi_registers.new_other\[9\] rbzero.spi_registers.spi_buffer\[9\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__mux2_1
X_20580_ _07685_ _07679_ _03451_ _03443_ rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__a32o_1
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19239_ rbzero.spi_registers.spi_done _02557_ _02558_ _02572_ vssd1 vssd1 vccd1 vccd1
+ _02771_ sky130_fd_sc_hd__and4b_1
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21201_ clknet_leaf_99_i_clk _00970_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21132_ clknet_leaf_94_i_clk _00901_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_21063_ net153 _00832_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20014_ _03259_ _03260_ net71 vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__o21ai_1
XFILLER_141_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ clknet_leaf_7_i_clk _00685_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_203_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20847_ clknet_leaf_49_i_clk _00616_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[3\]
+ sky130_fd_sc_hd__dfxtp_2
X_10600_ _03638_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11580_ _04357_ _04358_ _04329_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__mux2_1
XFILLER_195_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20778_ clknet_leaf_61_i_clk _00547_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
X_10531_ _03557_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__clkbuf_4
XFILLER_167_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ _05978_ _05982_ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__or3_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10462_ rbzero.tex_r0\[57\] rbzero.tex_r0\[56\] _03558_ vssd1 vssd1 vccd1 vccd1 _03566_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12201_ _04966_ net64 _04969_ _04970_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__a211o_1
X_13181_ _05844_ _05917_ _05834_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__a21o_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10393_ rbzero.tex_r1\[23\] rbzero.tex_r1\[24\] _03527_ vssd1 vssd1 vccd1 vccd1 _03528_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12132_ net9 net8 vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__nor2_2
XFILLER_151_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16940_ _09405_ _09444_ _09580_ vssd1 vssd1 vccd1 vccd1 _09581_ sky130_fd_sc_hd__a21o_1
XFILLER_2_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11014_ rbzero.tex_b0\[51\] rbzero.tex_b0\[50\] _03854_ vssd1 vssd1 vccd1 vccd1 _03856_
+ sky130_fd_sc_hd__mux2_1
X_16871_ _09510_ _09511_ vssd1 vssd1 vccd1 vccd1 _09512_ sky130_fd_sc_hd__nor2_1
XFILLER_42_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18610_ _02305_ _02306_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__xnor2_2
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _08440_ _08463_ vssd1 vssd1 vccd1 vccd1 _08467_ sky130_fd_sc_hd__nor2_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18541_ _10238_ _09434_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__nor2_1
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15753_ _08373_ _08390_ vssd1 vssd1 vccd1 vccd1 _08398_ sky130_fd_sc_hd__and2b_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _05673_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__buf_2
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ _05741_ _07383_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__or2_1
X_11916_ _04329_ _04691_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__or2_1
X_18472_ _09661_ _09611_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__and2_1
X_15684_ _08328_ vssd1 vssd1 vccd1 vccd1 _08329_ sky130_fd_sc_hd__buf_4
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12896_ _05609_ _05619_ _05622_ _05566_ _05562_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__o311a_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _09434_ _09988_ vssd1 vssd1 vccd1 vccd1 _09990_ sky130_fd_sc_hd__and2_1
X_14635_ _05931_ _07371_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__or2_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ rbzero.tex_g1\[37\] rbzero.tex_g1\[36\] _04392_ vssd1 vssd1 vccd1 vccd1 _04624_
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _09679_ _09659_ vssd1 vssd1 vccd1 vccd1 _09921_ sky130_fd_sc_hd__or2b_1
XFILLER_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14566_ _07294_ _07301_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__nor2_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _04140_ _04539_ _04555_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__or3_1
XFILLER_186_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13517_ _06206_ _06200_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__or2b_1
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16305_ _08945_ vssd1 vssd1 vccd1 vccd1 _08950_ sky130_fd_sc_hd__inv_2
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10729_ _03557_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__clkbuf_4
X_17285_ _09854_ _09855_ _09856_ vssd1 vssd1 vccd1 vccd1 _09858_ sky130_fd_sc_hd__o21a_1
X_14497_ _07184_ _07193_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16236_ _08825_ _08880_ vssd1 vssd1 vccd1 vccd1 _08881_ sky130_fd_sc_hd__xor2_1
X_19024_ _02643_ vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13448_ _06183_ _06184_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__and2_1
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16167_ _08794_ _08796_ vssd1 vssd1 vccd1 vccd1 _08812_ sky130_fd_sc_hd__xnor2_1
X_13379_ _05979_ _05909_ _05920_ _05900_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__or4b_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15118_ _04462_ rbzero.debug_overlay.vplaneX\[-7\] _07774_ _07775_ vssd1 vssd1 vccd1
+ vccd1 _07776_ sky130_fd_sc_hd__o22a_1
XFILLER_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16098_ _08722_ _08721_ vssd1 vssd1 vccd1 vccd1 _08743_ sky130_fd_sc_hd__xor2_1
XFILLER_5_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15049_ _07710_ _07711_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__or2b_1
X_19926_ rbzero.debug_overlay.playerY\[1\] _03193_ _03222_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _00999_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_74_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19857_ rbzero.pov.ready_buffer\[68\] _03164_ _03155_ _03169_ vssd1 vssd1 vccd1 vccd1
+ _03170_ sky130_fd_sc_hd__o211a_1
XFILLER_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18808_ _05204_ _02488_ _02489_ _10173_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__a31o_1
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19788_ rbzero.pov.spi_buffer\[67\] rbzero.pov.spi_buffer\[68\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03123_ sky130_fd_sc_hd__mux2_1
XFILLER_110_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_89_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18739_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.stepDistY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__nand2_1
XFILLER_3_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20701_ clknet_leaf_51_i_clk _00485_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_180_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20632_ clknet_leaf_12_i_clk _00416_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20563_ rbzero.traced_texVinit\[6\] _03443_ _09771_ _09597_ vssd1 vssd1 vccd1 vccd1
+ _01414_ sky130_fd_sc_hd__a22o_1
XFILLER_177_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20494_ _03389_ _03390_ _03391_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__and3_1
XFILLER_180_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20251__270 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__inv_2
XFILLER_191_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21115_ net205 _00884_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21046_ clknet_leaf_76_i_clk _00815_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ rbzero.map_rom.f4 _05497_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__or2_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _04470_ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__and2_1
XFILLER_91_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12681_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__nand2_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _07144_ _07156_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__xor2_1
XFILLER_187_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11632_ _04206_ _04374_ _04410_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__and3b_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14351_ _07006_ _07026_ _07087_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__a21oi_1
X_11563_ _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__buf_6
XFILLER_196_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13302_ _06022_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__xnor2_1
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10514_ _03593_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__clkbuf_1
X_17070_ _09560_ _09561_ vssd1 vssd1 vccd1 vccd1 _09710_ sky130_fd_sc_hd__nand2_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14282_ _06774_ _07018_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__nand2_1
XFILLER_183_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11494_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _04273_ vssd1 vssd1 vccd1 vccd1 _04274_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20334__345 clknet_1_1__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__inv_2
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16021_ _08621_ _08665_ vssd1 vssd1 vccd1 vccd1 _08666_ sky130_fd_sc_hd__xnor2_2
X_13233_ _05951_ _05924_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__nand2_1
X_10445_ _03474_ _03554_ _03555_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__or3_2
XFILLER_100_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13164_ _05743_ _05754_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__and2_2
X_10376_ rbzero.tex_r1\[31\] rbzero.tex_r1\[32\] _03516_ vssd1 vssd1 vccd1 vccd1 _03519_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12115_ gpout0.vpos\[7\] vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__buf_2
XFILLER_152_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17972_ _01670_ _01673_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__and2_1
XFILLER_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13095_ _05740_ _05831_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__nand2_1
XFILLER_3_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19711_ rbzero.pov.spi_buffer\[30\] rbzero.pov.spi_buffer\[31\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03083_ sky130_fd_sc_hd__mux2_1
X_12046_ _04318_ _04810_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nor2_1
XFILLER_172_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16923_ _07585_ _09431_ _09563_ _09085_ vssd1 vssd1 vccd1 vccd1 _09564_ sky130_fd_sc_hd__a211o_1
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03311_ _03311_ vssd1 vssd1 vccd1 vccd1 clknet_0__03311_ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16854_ _09492_ _09494_ vssd1 vssd1 vccd1 vccd1 _09495_ sky130_fd_sc_hd__nor2_1
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _07976_ _08215_ _08446_ _08449_ vssd1 vssd1 vccd1 vccd1 _08450_ sky130_fd_sc_hd__o31a_1
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16785_ _07598_ _09283_ _05209_ _09287_ vssd1 vssd1 vccd1 vccd1 _09427_ sky130_fd_sc_hd__or4_1
X_13997_ _06732_ _06733_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__or2_1
XFILLER_19_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20405__6 clknet_1_1__leaf__03037_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__inv_2
X_20380__387 clknet_1_1__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__inv_2
XFILLER_34_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18524_ _02138_ _02120_ _02221_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a21o_2
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12948_ _05577_ _05579_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__nand2_2
X_15736_ _08259_ _08238_ _08379_ _08380_ vssd1 vssd1 vccd1 vccd1 _08381_ sky130_fd_sc_hd__o31a_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18455_ _02151_ _02152_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__xor2_1
XFILLER_179_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15667_ _08306_ _08310_ _08311_ vssd1 vssd1 vccd1 vccd1 _08312_ sky130_fd_sc_hd__a21oi_1
X_12879_ _04030_ _05362_ _05363_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__and3_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ _09540_ vssd1 vssd1 vccd1 vccd1 _09973_ sky130_fd_sc_hd__clkbuf_4
XFILLER_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14618_ _07308_ _07315_ _07304_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__a21oi_1
X_18386_ _01982_ _01983_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__nand2_1
X_15598_ _08210_ _08213_ _07598_ _08002_ _05208_ vssd1 vssd1 vccd1 vccd1 _08243_ sky130_fd_sc_hd__a2111o_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17337_ _09605_ _09606_ _09734_ vssd1 vssd1 vccd1 vccd1 _09904_ sky130_fd_sc_hd__or3_1
X_14549_ _07270_ _07268_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__xor2_1
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17268_ _05531_ _09068_ vssd1 vssd1 vccd1 vccd1 _09843_ sky130_fd_sc_hd__nand2_1
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19007_ _02634_ vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__clkbuf_1
X_16219_ _08854_ _08861_ _08863_ vssd1 vssd1 vccd1 vccd1 _08864_ sky130_fd_sc_hd__a21oi_1
X_17199_ rbzero.wall_tracer.mapX\[7\] _05512_ vssd1 vssd1 vccd1 vccd1 _09783_ sky130_fd_sc_hd__and2_1
XFILLER_155_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19909_ _08070_ _03141_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__nor2_1
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21664_ clknet_leaf_34_i_clk _01433_ vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__03300_ clknet_0__03300_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03300_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20615_ clknet_leaf_71_i_clk _00011_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rcp_sel\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21595_ net136 _01364_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20546_ rbzero.traced_texa\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _03436_
+ sky130_fd_sc_hd__nand2_1
XFILLER_126_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20477_ rbzero.traced_texa\[-1\] rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1 _03378_
+ sky130_fd_sc_hd__or2_1
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20059__97 clknet_1_0__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__inv_2
XFILLER_121_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19606__60 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__inv_2
XFILLER_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13920_ _06598_ _06643_ _06653_ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__o211a_1
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21029_ clknet_leaf_13_i_clk _00798_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13851_ _06586_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__nand2_1
XFILLER_207_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19621__74 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__inv_2
XFILLER_76_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12802_ _05539_ _05543_ _05540_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__o21bai_1
XFILLER_28_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16570_ rbzero.wall_tracer.visualWallDist\[7\] _04015_ _08416_ _09211_ vssd1 vssd1
+ vccd1 vccd1 _09213_ sky130_fd_sc_hd__a31o_1
X_13782_ _06515_ _06518_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__or2_1
X_10994_ _03845_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_90_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15521_ _08155_ _08156_ _08164_ vssd1 vssd1 vccd1 vccd1 _08166_ sky130_fd_sc_hd__nor3_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _05424_ _05480_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__xnor2_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18240_ _10094_ _09162_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__nor2_1
XFILLER_163_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15452_ _08096_ vssd1 vssd1 vccd1 vccd1 _08097_ sky130_fd_sc_hd__clkbuf_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _05411_ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__nor2_8
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14403_ _07136_ _07137_ _07139_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__a21oi_1
XFILLER_169_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11615_ rbzero.tex_r1\[41\] rbzero.tex_r1\[40\] _04392_ vssd1 vssd1 vccd1 vccd1 _04394_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18171_ _10248_ _09973_ _01746_ _01871_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__o31a_1
XFILLER_129_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15383_ rbzero.debug_overlay.playerX\[-1\] rbzero.debug_overlay.playerX\[-2\] _08027_
+ vssd1 vssd1 vccd1 vccd1 _08028_ sky130_fd_sc_hd__or3_4
XFILLER_169_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12595_ _05347_ _05348_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__and2_1
XFILLER_196_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17122_ _04430_ _09750_ vssd1 vssd1 vccd1 vccd1 _09756_ sky130_fd_sc_hd__and2_1
X_14334_ _06705_ _07060_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__xor2_1
X_11546_ _04325_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__inv_2
XFILLER_11_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17053_ _09555_ vssd1 vssd1 vccd1 vccd1 _09693_ sky130_fd_sc_hd__buf_4
XFILLER_167_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14265_ _06999_ _07000_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__and2_1
X_11477_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _04213_ vssd1 vssd1 vccd1 vccd1 _04257_
+ sky130_fd_sc_hd__mux2_1
X_16004_ _08641_ _08647_ vssd1 vssd1 vccd1 vccd1 _08649_ sky130_fd_sc_hd__nor2_1
X_13216_ _05725_ _05723_ _05893_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__mux2_1
X_10428_ rbzero.tex_r1\[6\] rbzero.tex_r1\[7\] _03538_ vssd1 vssd1 vccd1 vccd1 _03546_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14196_ _06805_ _06668_ _06928_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__o21bai_1
XFILLER_48_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _05820_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__clkbuf_4
X_10359_ rbzero.tex_r1\[39\] net54 _03505_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__mux2_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17955_ _01492_ _01538_ _01657_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__a21oi_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _05640_ _05645_ _05648_ _05687_ _05795_ _05801_ vssd1 vssd1 vccd1 vccd1 _05815_
+ sky130_fd_sc_hd__mux4_1
XFILLER_140_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _09542_ _09423_ _09546_ vssd1 vssd1 vccd1 vccd1 _09547_ sky130_fd_sc_hd__o21a_1
X_12029_ _04244_ _04795_ _04803_ _04116_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a31o_1
XFILLER_65_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17886_ _01586_ _01587_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__and2_1
XFILLER_120_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16837_ _09403_ _09386_ vssd1 vssd1 vccd1 vccd1 _09478_ sky130_fd_sc_hd__or2b_1
XFILLER_81_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19556_ rbzero.pov.spi_counter\[2\] _03022_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__and2_1
X_16768_ _08284_ _09126_ _09276_ _08283_ vssd1 vssd1 vccd1 vccd1 _09410_ sky130_fd_sc_hd__o22a_1
XFILLER_94_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18507_ _02099_ _02065_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__or2b_1
XFILLER_20_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15719_ _08338_ _08339_ _08343_ vssd1 vssd1 vccd1 vccd1 _08364_ sky130_fd_sc_hd__o21ba_1
X_19487_ _02965_ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__xnor2_1
X_16699_ _09207_ _09330_ _09328_ vssd1 vssd1 vccd1 vccd1 _09341_ sky130_fd_sc_hd__a21bo_1
XFILLER_181_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18438_ _02135_ _02136_ _09780_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18369_ _02066_ _02067_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__nor2_1
XFILLER_187_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21380_ net301 _01149_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20363__371 clknet_1_0__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__inv_2
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21647_ clknet_leaf_32_i_clk _01416_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11400_ rbzero.row_render.size\[9\] _04153_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__nor2_1
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12380_ _04867_ _05145_ _05146_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__and3_1
XFILLER_197_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21578_ net499 _01347_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_70 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ rbzero.traced_texVinit\[11\] rbzero.texV\[11\] vssd1 vssd1 vccd1 vccd1 _04111_
+ sky130_fd_sc_hd__xor2_1
XFILLER_10_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20529_ _03416_ _03419_ _03417_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14050_ _06773_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__inv_2
XFILLER_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11262_ _04040_ _04041_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__nand2_2
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13001_ _05733_ _05735_ _05736_ _05737_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__a211o_1
XFILLER_107_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11193_ _03942_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__inv_2
XFILLER_95_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17740_ _10232_ _10197_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__or2b_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14952_ _04019_ _07643_ _07644_ _07642_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__o211a_1
XFILLER_43_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13903_ _06616_ _06639_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__xnor2_2
XFILLER_43_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17671_ _10112_ _10120_ _10119_ vssd1 vssd1 vccd1 vccd1 _10236_ sky130_fd_sc_hd__a21oi_2
X_14883_ rbzero.wall_tracer.visualWallDist\[-12\] _07595_ vssd1 vssd1 vccd1 vccd1
+ _07596_ sky130_fd_sc_hd__or2_1
XFILLER_47_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19410_ _02878_ _02880_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__or2b_1
X_16622_ _09263_ _09264_ vssd1 vssd1 vccd1 vccd1 _09265_ sky130_fd_sc_hd__nand2_1
X_13834_ _06569_ _06570_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__nand2_1
XFILLER_62_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19341_ _02830_ _02831_ _02829_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__nand3b_1
XFILLER_188_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ _06065_ _06031_ _06002_ _05877_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__a2bb2o_1
X_16553_ _09194_ _09196_ vssd1 vssd1 vccd1 vccd1 _09197_ sky130_fd_sc_hd__nor2_1
X_10977_ _03836_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15504_ rbzero.wall_tracer.visualWallDist\[3\] _08148_ vssd1 vssd1 vccd1 vccd1 _08149_
+ sky130_fd_sc_hd__nand2_4
XFILLER_206_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12716_ _05437_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__inv_2
X_19272_ _02783_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__inv_2
XFILLER_188_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16484_ _08180_ _08971_ vssd1 vssd1 vccd1 vccd1 _09128_ sky130_fd_sc_hd__nor2_1
X_13696_ _06383_ _06432_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__nand2_1
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18223_ _01833_ _01836_ _01921_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__nand3_1
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15435_ rbzero.debug_overlay.playerY\[-2\] _08029_ vssd1 vssd1 vccd1 vccd1 _08080_
+ sky130_fd_sc_hd__xor2_1
X_12647_ _03935_ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18154_ _01819_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__xnor2_1
X_15366_ _07997_ _08009_ _08010_ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12578_ _05288_ _05319_ _05323_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__o21ai_1
XFILLER_172_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20191__216 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__inv_2
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ _09470_ _09743_ _09600_ _09742_ vssd1 vssd1 vccd1 vccd1 _09745_ sky130_fd_sc_hd__a211o_1
XFILLER_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11529_ _04242_ _04298_ _04207_ _04308_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__o211a_1
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14317_ _07050_ _07052_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__and2_1
X_18085_ _01684_ _01685_ _01785_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__and3_1
XFILLER_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15297_ _07913_ _07924_ _07932_ _07941_ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__or4_1
XFILLER_116_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17036_ _08383_ _09674_ _09531_ _09675_ vssd1 vssd1 vccd1 vccd1 _09676_ sky130_fd_sc_hd__o31a_1
X_14248_ _06907_ _06908_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__or2_1
XFILLER_171_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14179_ _06905_ _06913_ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__or2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18987_ rbzero.pov.spi_buffer\[26\] rbzero.pov.ready_buffer\[26\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02624_ sky130_fd_sc_hd__mux2_1
XFILLER_61_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _01635_ _01639_ _01640_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__nand3_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17869_ _01448_ _01571_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20880_ clknet_leaf_98_i_clk _00649_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19600__55 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__inv_2
XFILLER_207_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19539_ rbzero.wall_tracer.rayAddendY\[10\] rbzero.wall_tracer.rayAddendY\[9\] _03001_
+ _02906_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__or4bb_1
XFILLER_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03039_ clknet_0__03039_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03039_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21501_ net422 _01270_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21432_ net353 _01201_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21363_ net284 _01132_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21294_ net215 _01063_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10900_ _03796_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__clkbuf_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11880_ rbzero.tex_g1\[31\] _04135_ _04136_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__and3_1
XFILLER_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_109 vssd1 vssd1 vccd1 vccd1 ones[3] top_ew_algofoogle_109/LO sky130_fd_sc_hd__conb_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10831_ rbzero.tex_g0\[10\] rbzero.tex_g0\[9\] _03751_ vssd1 vssd1 vccd1 vccd1 _03760_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13550_ _05990_ _05975_ _05984_ _05991_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__o22a_1
XFILLER_73_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10762_ rbzero.tex_g0\[43\] rbzero.tex_g0\[42\] _03718_ vssd1 vssd1 vccd1 vccd1 _03724_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12501_ _05254_ rbzero.wall_tracer.trackDistX\[2\] _05255_ rbzero.wall_tracer.trackDistX\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__o22a_1
X_13481_ _06214_ _06217_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__xnor2_1
X_10693_ _03687_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15220_ _07820_ rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 _07871_
+ sky130_fd_sc_hd__or2_1
XFILLER_139_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12432_ _04002_ _03914_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__nor2_1
XFILLER_148_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15151_ _07804_ _07806_ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__or2_1
X_12363_ _04883_ _04884_ _05083_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__mux2_1
XFILLER_5_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14102_ _06821_ _06837_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__nor2_1
X_11314_ _04065_ _04068_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__and2_1
XFILLER_181_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15082_ rbzero.debug_overlay.vplaneX\[0\] vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__buf_2
XFILLER_114_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12294_ net49 _05044_ _05046_ net52 vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__a22o_1
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14033_ _06615_ _06641_ _06642_ _06657_ _06769_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__a311oi_4
X_18910_ _02557_ _02573_ _02578_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__and3_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11245_ _04028_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__inv_2
XFILLER_106_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19890_ _03193_ _03195_ _03196_ _03157_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__o211a_1
XFILLER_84_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18841_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.stepDistY\[6\] vssd1
+ vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__and2_1
XFILLER_68_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11176_ _03960_ _03961_ _03962_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__and4_1
XFILLER_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18772_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.stepDistY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__nand2_1
X_15984_ _08559_ _08623_ _08624_ _08628_ vssd1 vssd1 vccd1 vccd1 _08629_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_76_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17723_ _10285_ _10287_ vssd1 vssd1 vccd1 vccd1 _10288_ sky130_fd_sc_hd__xor2_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14935_ rbzero.wall_tracer.visualWallDist\[3\] _07618_ vssd1 vssd1 vccd1 vccd1 _07633_
+ sky130_fd_sc_hd__or2_1
XFILLER_48_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17654_ _09522_ _08425_ _10218_ vssd1 vssd1 vccd1 vccd1 _10219_ sky130_fd_sc_hd__or3_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14866_ _05929_ _07456_ _07581_ _07487_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__o31a_2
XFILLER_35_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16605_ _09243_ _08059_ _09247_ vssd1 vssd1 vccd1 vccd1 _09248_ sky130_fd_sc_hd__or3_1
XFILLER_51_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13817_ _06376_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__xor2_1
XFILLER_63_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17585_ _10147_ _10150_ vssd1 vssd1 vccd1 vccd1 _10151_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14797_ _07473_ _07471_ _07526_ _07527_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__o211a_1
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19324_ _02818_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__clkbuf_1
X_16536_ _09178_ _09179_ vssd1 vssd1 vccd1 vccd1 _09180_ sky130_fd_sc_hd__and2_1
XFILLER_50_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13748_ _06383_ _06432_ _06484_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__a21oi_1
XFILLER_177_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19255_ _02780_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__clkbuf_1
XFILLER_149_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16467_ _09091_ _08968_ _09109_ vssd1 vssd1 vccd1 vccd1 _09111_ sky130_fd_sc_hd__and3_1
XFILLER_148_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13679_ _06395_ _06415_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18206_ _01905_ _01799_ _01801_ _05203_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__a31o_1
X_15418_ _08059_ _08062_ vssd1 vssd1 vccd1 vccd1 _08063_ sky130_fd_sc_hd__nor2_1
X_19186_ rbzero.spi_registers.new_leak\[4\] _02733_ vssd1 vssd1 vccd1 vccd1 _02738_
+ sky130_fd_sc_hd__or2_1
X_16398_ _09040_ _09042_ vssd1 vssd1 vccd1 vccd1 _09043_ sky130_fd_sc_hd__xnor2_1
XFILLER_191_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18137_ _01836_ _01837_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__and2_1
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15349_ _07925_ _07992_ _07993_ vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__a21oi_4
XFILLER_172_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18068_ _01753_ _01768_ _01769_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__nand3_1
XFILLER_160_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17019_ _09528_ _09535_ _09658_ vssd1 vssd1 vccd1 vccd1 _09659_ sky130_fd_sc_hd__a21o_1
X_20030_ _09753_ _03267_ _03271_ _03272_ _04883_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__a32o_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20932_ clknet_leaf_78_i_clk _00701_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20863_ clknet_leaf_0_i_clk _00632_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20794_ clknet_leaf_46_i_clk _00563_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20174__200 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__inv_2
XFILLER_10_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21415_ net336 _01184_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21346_ net267 _01115_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21277_ clknet_leaf_95_i_clk _01046_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[0\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11030_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _03854_ vssd1 vssd1 vccd1 vccd1 _03864_
+ sky130_fd_sc_hd__mux2_1
XFILLER_131_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12981_ _05598_ _05717_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__xor2_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _07431_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__inv_2
XFILLER_85_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11932_ _04210_ _04703_ _04707_ _04232_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a211o_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ rbzero.tex_g1\[3\] _04135_ _04136_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__and3_1
X_14651_ _07107_ _07356_ _07387_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__a21bo_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13602_ _05995_ _06113_ _06057_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__a21oi_2
XFILLER_14_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10814_ _03717_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__clkbuf_4
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _09926_ _09935_ vssd1 vssd1 vccd1 vccd1 _09937_ sky130_fd_sc_hd__or2_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _04254_ _04567_ _04571_ _04241_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a211o_1
X_14582_ _07294_ _07301_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__nand2_1
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16321_ _08964_ _08965_ vssd1 vssd1 vccd1 vccd1 _08966_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10745_ _03714_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__clkbuf_1
X_13533_ _06183_ _06222_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__nor2_1
XFILLER_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19040_ rbzero.pov.spi_buffer\[51\] rbzero.pov.ready_buffer\[51\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02652_ sky130_fd_sc_hd__mux2_1
X_16252_ _08893_ _08894_ _08896_ vssd1 vssd1 vccd1 vccd1 _08897_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13464_ _05923_ _05989_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__nand2_2
X_10676_ _03678_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12415_ _05146_ net66 _05181_ net36 vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__a211o_1
XFILLER_127_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15203_ _03913_ _07853_ _07854_ _07855_ rbzero.wall_tracer.rayAddendX\[7\] vssd1
+ vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__a32o_1
X_16183_ _08194_ _08491_ vssd1 vssd1 vccd1 vccd1 _08828_ sky130_fd_sc_hd__or2_1
X_13395_ _05824_ _06066_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__or2_1
XFILLER_51_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12346_ _05101_ _05111_ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__o21ba_1
XFILLER_182_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15134_ _07730_ rbzero.debug_overlay.vplaneX\[-5\] vssd1 vssd1 vccd1 vccd1 _07791_
+ sky130_fd_sc_hd__xor2_1
XFILLER_114_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15065_ rbzero.wall_tracer.rayAddendX\[-2\] _07726_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07727_ sky130_fd_sc_hd__mux2_1
X_19942_ rbzero.debug_overlay.playerY\[5\] vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__inv_2
X_12277_ _05032_ net20 vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__nor2_2
XFILLER_141_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14016_ _06680_ _06668_ _06714_ _06716_ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__o31ai_1
X_11228_ _04012_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__buf_4
XFILLER_141_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19873_ rbzero.debug_overlay.playerX\[3\] _03143_ _03182_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _00986_ sky130_fd_sc_hd__a211o_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18824_ rbzero.wall_tracer.trackDistY\[4\] rbzero.wall_tracer.stepDistY\[4\] vssd1
+ vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__nor2_1
X_11159_ rbzero.debug_overlay.playerX\[2\] _03929_ _03936_ rbzero.debug_overlay.playerX\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__o22a_1
XFILLER_191_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18755_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.stepDistY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__or2_1
X_15967_ _08586_ _08608_ vssd1 vssd1 vccd1 vccd1 _08612_ sky130_fd_sc_hd__nor2_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17706_ _10270_ vssd1 vssd1 vccd1 vccd1 _10271_ sky130_fd_sc_hd__buf_4
X_14918_ _04019_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__clkbuf_4
X_18686_ _02325_ _02381_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__xnor2_2
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ _08539_ _08541_ _08542_ vssd1 vssd1 vccd1 vccd1 _08543_ sky130_fd_sc_hd__a21oi_2
X_17637_ _09368_ _10200_ _10201_ vssd1 vssd1 vccd1 vccd1 _10202_ sky130_fd_sc_hd__o21bai_1
X_14849_ rbzero.wall_tracer.stepDistY\[5\] _07568_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07569_ sky130_fd_sc_hd__mux2_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17568_ _05211_ _09699_ _10128_ vssd1 vssd1 vccd1 vccd1 _10134_ sky130_fd_sc_hd__o21ai_2
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19307_ _02809_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__clkbuf_1
X_16519_ _05209_ _09162_ vssd1 vssd1 vccd1 vccd1 _09163_ sky130_fd_sc_hd__or2_1
XFILLER_143_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17499_ _10062_ _10063_ vssd1 vssd1 vccd1 vccd1 _10065_ sky130_fd_sc_hd__nand2_1
XFILLER_176_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19238_ rbzero.spi_registers.vshift\[5\] _02762_ _02770_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00763_ sky130_fd_sc_hd__o211a_1
XFILLER_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19169_ rbzero.spi_registers.got_new_vinf vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__inv_2
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21200_ clknet_leaf_99_i_clk _00969_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ss_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_117_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21131_ clknet_leaf_94_i_clk _00900_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21062_ net152 _00831_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20013_ _04883_ _04992_ _03257_ _04884_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__or4b_1
XFILLER_28_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20206__229 clknet_1_0__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__inv_2
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20915_ clknet_leaf_6_i_clk _00684_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20846_ clknet_leaf_49_i_clk _00615_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20777_ clknet_leaf_61_i_clk _00546_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10530_ _03601_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10461_ _03565_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__clkbuf_1
X_12200_ _04966_ _04738_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__nor2_1
X_13180_ _05842_ _05916_ _05807_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__mux2_1
XFILLER_202_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10392_ _03482_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__clkbuf_4
XFILLER_159_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12131_ net61 _04836_ _04839_ _04902_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__o31a_2
XFILLER_151_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21329_ net250 _01098_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12062_ clknet_opt_5_0_i_clk vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__buf_1
XFILLER_172_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11013_ _03855_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16870_ _09507_ _09509_ vssd1 vssd1 vccd1 vccd1 _09511_ sky130_fd_sc_hd__and2_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _08169_ _08465_ vssd1 vssd1 vccd1 vccd1 _08466_ sky130_fd_sc_hd__nor2_2
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18540_ _01737_ _10266_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__nor2_1
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _08392_ _08396_ vssd1 vssd1 vccd1 vccd1 _08397_ sky130_fd_sc_hd__xnor2_2
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _05638_ _05649_ _05687_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__or3_2
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _07106_ _07415_ _07416_ _07417_ _05742_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__o311ai_2
X_18471_ _02167_ _02168_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__xnor2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _04290_ vssd1 vssd1 vccd1 vccd1 _04691_
+ sky130_fd_sc_hd__mux2_1
X_20146__176 clknet_1_1__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__inv_2
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _08148_ _08037_ _08038_ vssd1 vssd1 vccd1 vccd1 _08328_ sky130_fd_sc_hd__a21oi_4
XFILLER_205_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _05623_ _05626_ _05628_ _05631_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__o211a_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _09434_ _09988_ vssd1 vssd1 vccd1 vccd1 _09989_ sky130_fd_sc_hd__nand2_1
XFILLER_166_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14634_ _07366_ _07370_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__nand2_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ rbzero.tex_g1\[39\] rbzero.tex_g1\[38\] _04392_ vssd1 vssd1 vccd1 vccd1 _04623_
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _09678_ _09660_ vssd1 vssd1 vccd1 vccd1 _09920_ sky130_fd_sc_hd__or2b_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _04142_ _04546_ _04554_ _04143_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__o211a_1
XFILLER_13_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14565_ _07294_ _07301_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__and2_1
XFILLER_186_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16304_ _08941_ _08811_ vssd1 vssd1 vccd1 vccd1 _08949_ sky130_fd_sc_hd__and2_1
XFILLER_202_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10728_ _03705_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__clkbuf_1
X_13516_ _06251_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__and2_1
XFILLER_207_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17284_ _09854_ _09855_ _09856_ vssd1 vssd1 vccd1 vccd1 _09857_ sky130_fd_sc_hd__nor3_1
XFILLER_140_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14496_ _07227_ _07231_ _07232_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__a21o_1
XFILLER_158_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19023_ rbzero.pov.spi_buffer\[43\] rbzero.pov.ready_buffer\[43\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02643_ sky130_fd_sc_hd__mux2_1
X_16235_ _08816_ _08821_ vssd1 vssd1 vccd1 vccd1 _08880_ sky130_fd_sc_hd__nor2_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10659_ rbzero.tex_g1\[27\] rbzero.tex_g1\[28\] _03669_ vssd1 vssd1 vccd1 vccd1 _03670_
+ sky130_fd_sc_hd__mux2_1
X_13447_ _06177_ _06178_ _06182_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_8_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13378_ _06045_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__inv_2
X_16166_ _08808_ _08810_ vssd1 vssd1 vccd1 vccd1 _08811_ sky130_fd_sc_hd__xor2_4
XFILLER_170_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15117_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.debug_overlay.vplaneX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__nor2_1
XFILLER_114_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12329_ _05090_ _05093_ _05094_ _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__and4_1
X_20311__324 clknet_1_0__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__inv_2
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16097_ _08700_ _08709_ vssd1 vssd1 vccd1 vccd1 _08742_ sky130_fd_sc_hd__xnor2_2
XFILLER_173_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15048_ _04462_ rbzero.wall_tracer.rayAddendX\[-3\] vssd1 vssd1 vccd1 vccd1 _07711_
+ sky130_fd_sc_hd__nand2_1
X_19925_ rbzero.pov.ready_buffer\[54\] _03164_ _03197_ _03221_ vssd1 vssd1 vccd1 vccd1
+ _03222_ sky130_fd_sc_hd__o211a_1
XFILLER_69_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19856_ rbzero.debug_overlay.playerX\[0\] _08028_ _03168_ vssd1 vssd1 vccd1 vccd1
+ _03169_ sky130_fd_sc_hd__a21o_1
XFILLER_122_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18807_ _02481_ _02483_ _02486_ _02487_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__o211ai_2
XFILLER_110_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19787_ _03122_ vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__clkbuf_1
X_16999_ _09501_ _09504_ _09503_ vssd1 vssd1 vccd1 vccd1 _09639_ sky130_fd_sc_hd__a21bo_1
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18738_ rbzero.wall_tracer.trackDistY\[-7\] rbzero.wall_tracer.stepDistY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__or2_1
X_20401__26 clknet_1_0__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__inv_2
XFILLER_37_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18669_ _02167_ _02255_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__nand2_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20700_ clknet_leaf_56_i_clk _00484_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_51_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20631_ clknet_leaf_14_i_clk _00415_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20562_ _07831_ _09458_ rbzero.traced_texVinit\[5\] _09762_ vssd1 vssd1 vccd1 vccd1
+ _01413_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_149_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20493_ _03389_ _03390_ _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a21o_1
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21114_ net204 _00883_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20286__301 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__inv_2
XFILLER_8_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21045_ clknet_leaf_81_i_clk _00814_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _04473_ _04478_ gpout0.vpos\[5\] gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1
+ _04479_ sky130_fd_sc_hd__o211a_1
X_12680_ _05424_ _05425_ _05426_ _05427_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__o211a_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _04207_ _04383_ _04391_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a31o_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ clknet_leaf_44_i_clk _00598_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11562_ _04128_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__buf_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14350_ _07023_ _07025_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__nor2_1
XFILLER_126_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10513_ rbzero.tex_r0\[33\] rbzero.tex_r0\[32\] _03591_ vssd1 vssd1 vccd1 vccd1 _03593_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13301_ _06024_ _06029_ _06037_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__o21ai_2
XFILLER_13_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14281_ _06805_ _06761_ _06772_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__o21ai_1
X_11493_ _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__buf_4
XFILLER_171_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13232_ _05901_ _05904_ _05964_ _05968_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__a211o_1
X_16020_ _08654_ _08663_ _08664_ vssd1 vssd1 vccd1 vccd1 _08665_ sky130_fd_sc_hd__a21oi_1
XFILLER_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10444_ _03479_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__inv_12
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ _05846_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__nor2_1
X_10375_ _03518_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12114_ gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__buf_2
X_17971_ _01669_ _01670_ _01673_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__and3_1
X_13094_ _05829_ _05830_ _05778_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__mux2_1
XFILLER_152_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19710_ _03082_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__clkbuf_1
X_12045_ _04809_ _04810_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__xnor2_1
X_16922_ _07575_ _08983_ _09430_ _07586_ vssd1 vssd1 vccd1 vccd1 _09563_ sky130_fd_sc_hd__o31a_1
XFILLER_46_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03310_ _03310_ vssd1 vssd1 vccd1 vccd1 clknet_0__03310_ sky130_fd_sc_hd__clkbuf_16
XFILLER_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16853_ _08335_ _09165_ _09354_ _09493_ vssd1 vssd1 vccd1 vccd1 _09494_ sky130_fd_sc_hd__o31a_1
XFILLER_78_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15804_ _08202_ _08238_ _08448_ vssd1 vssd1 vccd1 vccd1 _08449_ sky130_fd_sc_hd__or3_1
XFILLER_20_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16784_ _08377_ _09138_ vssd1 vssd1 vccd1 vccd1 _09426_ sky130_fd_sc_hd__nor2_1
XFILLER_168_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13996_ _06731_ _06700_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__and2_1
XFILLER_206_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18523_ _02218_ _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__xnor2_2
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15735_ _08303_ _08378_ vssd1 vssd1 vccd1 vccd1 _08380_ sky130_fd_sc_hd__nand2_1
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12947_ _05673_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__or2_2
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _10248_ _10266_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__nor2_1
X_15666_ _08299_ _08305_ vssd1 vssd1 vccd1 vccd1 _08311_ sky130_fd_sc_hd__nor2_1
XFILLER_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12878_ _05561_ _05466_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__o21a_2
XFILLER_61_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17405_ _09957_ _09971_ vssd1 vssd1 vccd1 vccd1 _09972_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _07304_ _07308_ _07315_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__and3_1
X_18385_ _01955_ _01957_ _01954_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__a21bo_1
X_11829_ rbzero.tex_g1\[56\] _04272_ _04139_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__a21o_1
X_15597_ _08217_ _08225_ _05198_ vssd1 vssd1 vccd1 vccd1 _08242_ sky130_fd_sc_hd__o21ai_4
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17336_ rbzero.wall_tracer.trackDistX\[-1\] _09817_ _09897_ _09903_ vssd1 vssd1 vccd1
+ vccd1 _00588_ sky130_fd_sc_hd__o22a_1
XFILLER_144_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14548_ _07250_ _07272_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__xor2_1
XFILLER_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17267_ _09838_ _09839_ _09840_ vssd1 vssd1 vccd1 vccd1 _09842_ sky130_fd_sc_hd__o21a_1
XFILLER_174_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14479_ _07200_ _07215_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__and2_1
XFILLER_162_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19006_ rbzero.pov.spi_buffer\[35\] rbzero.pov.ready_buffer\[35\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02634_ sky130_fd_sc_hd__mux2_1
X_16218_ _08250_ _08331_ _08862_ vssd1 vssd1 vccd1 vccd1 _08863_ sky130_fd_sc_hd__and3_1
XFILLER_128_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17198_ rbzero.wall_tracer.mapX\[6\] _05512_ _09778_ vssd1 vssd1 vccd1 vccd1 _09782_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16149_ _08776_ _08793_ vssd1 vssd1 vccd1 vccd1 _08794_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19908_ rbzero.debug_overlay.playerY\[-4\] _03198_ _03208_ _03209_ vssd1 vssd1 vccd1
+ vccd1 _00994_ sky130_fd_sc_hd__o211a_1
XFILLER_130_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19839_ _05190_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__clkbuf_4
XFILLER_83_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20129__160 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__inv_2
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20281__297 clknet_1_0__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__inv_2
XFILLER_36_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21663_ clknet_leaf_34_i_clk _01432_ vssd1 vssd1 vccd1 vccd1 gpout2.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20614_ _03472_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21594_ net135 _01363_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20545_ rbzero.traced_texa\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _03435_
+ sky130_fd_sc_hd__or2_1
XFILLER_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20476_ _03374_ _03375_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__nor2_1
XFILLER_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21028_ clknet_leaf_11_i_clk _00797_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13850_ _06574_ _06585_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__or2_1
XFILLER_142_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12801_ rbzero.wall_tracer.mapY\[7\] _05404_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__nor2_1
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10993_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _03843_ vssd1 vssd1 vccd1 vccd1 _03845_
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13781_ _06503_ _06516_ _06517_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__and3_1
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15520_ _08155_ _08156_ _08164_ vssd1 vssd1 vccd1 vccd1 _08165_ sky130_fd_sc_hd__o21a_1
XFILLER_128_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20340__350 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__inv_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _05479_ _05425_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__nor2_2
XFILLER_163_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15451_ _07945_ _08091_ _08095_ vssd1 vssd1 vccd1 vccd1 _08096_ sky130_fd_sc_hd__o21ai_4
XFILLER_188_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ rbzero.wall_tracer.state\[1\] _05211_ _04017_ _05278_ _05281_ vssd1 vssd1
+ vccd1 vccd1 _05412_ sky130_fd_sc_hd__o221ai_4
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_73_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14402_ _06724_ _06663_ _07138_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__nor3_1
X_18170_ _01744_ _01745_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__nand2_1
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11614_ rbzero.tex_r1\[43\] rbzero.tex_r1\[42\] _04392_ vssd1 vssd1 vccd1 vccd1 _04393_
+ sky130_fd_sc_hd__mux2_1
X_15382_ rbzero.debug_overlay.playerX\[-3\] _07946_ vssd1 vssd1 vccd1 vccd1 _08027_
+ sky130_fd_sc_hd__or2_1
XFILLER_169_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12594_ _05289_ _05295_ _05303_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__a21o_1
X_17121_ _04426_ _09748_ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__nor2_1
X_20258__277 clknet_1_0__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__inv_2
X_14333_ _07067_ _07069_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__xor2_1
X_11545_ _04047_ _04311_ _04313_ _04324_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__a31o_4
XFILLER_204_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17052_ _09682_ _09691_ vssd1 vssd1 vccd1 vccd1 _09692_ sky130_fd_sc_hd__xnor2_4
X_11476_ _04210_ _04248_ _04255_ _04232_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__a211o_1
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14264_ _06999_ _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__nor2_1
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_88_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16003_ _08641_ _08647_ vssd1 vssd1 vccd1 vccd1 _08648_ sky130_fd_sc_hd__xor2_1
X_10427_ _03545_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__clkbuf_1
X_13215_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__clkbuf_4
X_14195_ _06923_ _06931_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ _03509_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__clkbuf_1
X_13146_ _05844_ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__nor2_1
XFILLER_97_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_11_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17954_ _01535_ _01537_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__nor2_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _05813_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__clkbuf_4
X_16905_ _09544_ _09545_ vssd1 vssd1 vccd1 vccd1 _09546_ sky130_fd_sc_hd__xnor2_1
X_12028_ _04797_ _04799_ _04802_ _04306_ _04241_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a221o_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17885_ _01586_ _01587_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__nor2_1
XFILLER_65_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16836_ _09362_ _09377_ _09375_ vssd1 vssd1 vccd1 vccd1 _09477_ sky130_fd_sc_hd__a21o_1
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19555_ _03027_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16767_ _08284_ _09276_ vssd1 vssd1 vccd1 vccd1 _09409_ sky130_fd_sc_hd__nor2_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13979_ _06245_ _06678_ _06715_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__or3b_1
XFILLER_80_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18506_ _02202_ _02203_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__nor2_1
XFILLER_207_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15718_ _08361_ _08362_ vssd1 vssd1 vccd1 vccd1 _08363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19486_ _02938_ _02956_ _02958_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__a21o_1
XFILLER_181_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16698_ _05194_ _09339_ _09340_ _07642_ vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__o211a_1
XFILLER_55_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18437_ _02132_ _02133_ _02134_ _05204_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__o31a_1
X_15649_ _08292_ _08293_ vssd1 vssd1 vccd1 vccd1 _08294_ sky130_fd_sc_hd__xnor2_2
XFILLER_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18368_ _01474_ _09350_ _01934_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__o21a_1
XFILLER_187_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17319_ _05532_ _09597_ vssd1 vssd1 vccd1 vccd1 _09888_ sky130_fd_sc_hd__and2_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18299_ _01885_ _01887_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__and2_1
XFILLER_186_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21646_ clknet_leaf_32_i_clk _01415_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21577_ net498 _01346_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_60 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_71 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _04048_ _04051_ _04109_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__o21ai_1
XANTENNA_82 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20528_ rbzero.traced_texa\[7\] rbzero.texV\[7\] vssd1 vssd1 vccd1 vccd1 _03421_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_153_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11261_ gpout0.vpos\[5\] gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__nor2_2
X_20459_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 _03363_
+ sky130_fd_sc_hd__and2_1
X_13000_ _05649_ _05695_ _05673_ _05696_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__or4_4
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11192_ _03933_ rbzero.map_rom.a6 rbzero.map_rom.i_row\[4\] _03974_ _03924_ vssd1
+ vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__o32a_1
XFILLER_133_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14951_ rbzero.wall_tracer.visualWallDist\[8\] _07594_ vssd1 vssd1 vccd1 vccd1 _07644_
+ sky130_fd_sc_hd__or2_1
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13902_ _06617_ _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__xor2_2
X_17670_ _10098_ _10106_ _10234_ vssd1 vssd1 vccd1 vccd1 _10235_ sky130_fd_sc_hd__a21o_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14882_ _07594_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__clkbuf_4
XFILLER_75_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16621_ _09241_ _09242_ _09262_ vssd1 vssd1 vccd1 vccd1 _09264_ sky130_fd_sc_hd__nand3_1
X_13833_ _05974_ _06245_ _06161_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__o21ai_1
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19340_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__or2_1
X_16552_ rbzero.debug_overlay.playerX\[-5\] _07971_ _09195_ vssd1 vssd1 vccd1 vccd1
+ _09196_ sky130_fd_sc_hd__o21ai_2
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13764_ _06065_ _05947_ _05975_ _05984_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__or4_1
X_10976_ rbzero.tex_b1\[4\] rbzero.tex_b1\[5\] _03828_ vssd1 vssd1 vccd1 vccd1 _03836_
+ sky130_fd_sc_hd__mux2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15503_ _04014_ vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__buf_6
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12715_ _05462_ _05440_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__nand2_1
X_19271_ _02789_ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__clkbuf_1
X_16483_ _09126_ _08194_ vssd1 vssd1 vccd1 vccd1 _09127_ sky130_fd_sc_hd__nor2_1
XFILLER_206_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13695_ _05824_ _06240_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__nor2_1
X_18222_ _01833_ _01836_ _01921_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__a21o_1
XFILLER_70_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15434_ _08077_ _08078_ _05496_ vssd1 vssd1 vccd1 vccd1 _08079_ sky130_fd_sc_hd__mux2_1
X_12646_ _05374_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__clkbuf_4
XFILLER_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18153_ _01821_ _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15365_ _07977_ _07995_ _07981_ _07989_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__or4_1
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12577_ _05329_ _05330_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__nand2_1
XFILLER_8_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17104_ _09461_ _09465_ _09600_ _09742_ _09743_ vssd1 vssd1 vccd1 vccd1 _09744_ sky130_fd_sc_hd__o311a_1
XFILLER_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _07050_ _07052_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__nor2_1
X_18084_ _01684_ _01685_ _01785_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__a21oi_1
X_11528_ _04230_ _04301_ _04232_ _04307_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__a211o_1
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15296_ _07940_ vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__clkbuf_4
XFILLER_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17035_ _09396_ _09669_ vssd1 vssd1 vccd1 vccd1 _09675_ sky130_fd_sc_hd__nand2_1
X_14247_ _06981_ _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__and2_1
X_11459_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _04214_ vssd1 vssd1 vccd1 vccd1 _04239_
+ sky130_fd_sc_hd__mux2_1
XFILLER_113_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14178_ _06885_ _06911_ _06914_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__and3_1
XFILLER_180_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13129_ _05715_ _05721_ _05734_ _05718_ _05777_ _05801_ vssd1 vssd1 vccd1 vccd1 _05866_
+ sky130_fd_sc_hd__mux4_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _02623_ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__clkbuf_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17937_ _01636_ _01637_ _01638_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__a21o_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17868_ _01569_ _01570_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__nor2_1
XFILLER_66_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19597__52 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__inv_2
XFILLER_4_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16819_ _09458_ _09460_ vssd1 vssd1 vccd1 vccd1 _09461_ sky130_fd_sc_hd__nor2_1
X_17799_ _09668_ _09973_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__nor2_1
XFILLER_4_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19538_ _03009_ _03013_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__nand2_1
XFILLER_50_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03038_ clknet_0__03038_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03038_
+ sky130_fd_sc_hd__clkbuf_16
X_19469_ _02948_ _02949_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__nand2_1
XFILLER_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21500_ net421 _01269_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21431_ net352 _01200_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21362_ net283 _01131_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21293_ net214 _01062_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10830_ _03759_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _03723_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ rbzero.wall_tracer.trackDistY\[1\] vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__inv_2
XFILLER_198_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10692_ rbzero.tex_g1\[11\] rbzero.tex_g1\[12\] _03680_ vssd1 vssd1 vccd1 vccd1 _03687_
+ sky130_fd_sc_hd__mux2_1
XFILLER_125_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13480_ _05921_ _06176_ _06215_ _06216_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__a31oi_1
XFILLER_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12431_ _05192_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21629_ clknet_leaf_46_i_clk _01398_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15150_ _07792_ _07791_ _07805_ _07775_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__o22a_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12362_ _05124_ _05129_ _05081_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__o21a_2
XFILLER_148_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14101_ _06821_ _06837_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__xor2_1
XFILLER_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11313_ _04081_ _04089_ _04092_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__o21a_1
X_12293_ _05055_ net22 vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__nand2_1
X_15081_ _07729_ _07733_ _07731_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__a21bo_1
XFILLER_180_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14032_ _06016_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__clkbuf_4
X_11244_ _03912_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__nor2_2
XFILLER_141_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18840_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.stepDistY\[6\] vssd1
+ vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__nor2_1
X_11175_ rbzero.otherx\[3\] _03936_ _03921_ rbzero.othery\[3\] _03963_ vssd1 vssd1
+ vccd1 vccd1 _03964_ sky130_fd_sc_hd__o221a_1
XFILLER_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20069__106 clknet_1_0__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__inv_2
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18771_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.stepDistY\[-3\] vssd1
+ vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__or2_1
XFILLER_110_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15983_ _08625_ _08627_ vssd1 vssd1 vccd1 vccd1 _08628_ sky130_fd_sc_hd__xnor2_1
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17722_ _10048_ _10159_ _10286_ vssd1 vssd1 vccd1 vccd1 _10287_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14934_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.trackDistX\[3\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__mux2_1
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17653_ _10074_ _10217_ vssd1 vssd1 vccd1 vccd1 _10218_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14865_ _07435_ _07436_ _07433_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16604_ _09244_ _09246_ vssd1 vssd1 vccd1 vccd1 _09247_ sky130_fd_sc_hd__nand2_1
X_13816_ _06336_ _06375_ _06424_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__o21ba_1
XFILLER_35_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17584_ _10148_ _10149_ _10005_ _10006_ _09986_ vssd1 vssd1 vccd1 vccd1 _10150_ sky130_fd_sc_hd__a32o_2
XFILLER_17_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14796_ _05834_ _05800_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__nor2_2
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19323_ rbzero.spi_registers.new_vshift\[4\] rbzero.spi_registers.spi_buffer\[4\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__mux2_1
X_16535_ _09161_ _09166_ _09177_ vssd1 vssd1 vccd1 vccd1 _09179_ sky130_fd_sc_hd__o21bai_1
XFILLER_32_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13747_ _06065_ _06240_ _06161_ _05824_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__o22a_1
XFILLER_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10959_ rbzero.tex_b1\[12\] rbzero.tex_b1\[13\] _03817_ vssd1 vssd1 vccd1 vccd1 _03827_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19254_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_sky\[5\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__mux2_1
XFILLER_149_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16466_ _09091_ _08968_ _09109_ vssd1 vssd1 vccd1 vccd1 _09110_ sky130_fd_sc_hd__a21oi_1
X_13678_ _06396_ _06413_ _06414_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18205_ _01799_ _01801_ _01905_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15417_ _05193_ _07465_ _08061_ vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__a21oi_4
X_19185_ rbzero.floor_leak\[3\] _02732_ _02737_ _02722_ vssd1 vssd1 vccd1 vccd1 _00743_
+ sky130_fd_sc_hd__o211a_1
X_12629_ _03933_ _05374_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__nor2_1
X_16397_ _08430_ _09041_ vssd1 vssd1 vccd1 vccd1 _09042_ sky130_fd_sc_hd__nor2_1
XFILLER_106_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18136_ _01826_ _01835_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__or2_1
XFILLER_185_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15348_ _07904_ rbzero.wall_tracer.stepDistY\[-3\] _05206_ vssd1 vssd1 vccd1 vccd1
+ _07993_ sky130_fd_sc_hd__a21o_1
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18067_ _01766_ _01767_ _01754_ _01647_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__o211ai_2
XFILLER_176_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15279_ _07923_ vssd1 vssd1 vccd1 vccd1 _07924_ sky130_fd_sc_hd__buf_2
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17018_ _09533_ _09534_ vssd1 vssd1 vccd1 vccd1 _09658_ sky130_fd_sc_hd__nor2_1
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _02614_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__clkbuf_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20931_ clknet_leaf_77_i_clk _00700_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20862_ clknet_leaf_0_i_clk _00631_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20793_ clknet_leaf_28_i_clk _00562_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21414_ net335 _01183_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21345_ net266 _01114_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21276_ clknet_leaf_93_i_clk _01045_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-1\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_150_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20227_ clknet_1_1__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__buf_1
XFILLER_1_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12980_ _05594_ _05596_ _05628_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__o21a_1
XFILLER_76_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _04704_ _04705_ _04706_ _04219_ _04254_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__o221a_1
XFILLER_17_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19576__33 clknet_1_1__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__inv_2
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14650_ _05793_ _07369_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__nand2_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _04637_ _04638_ _04224_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__mux2_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _05988_ _06337_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__xnor2_1
XFILLER_72_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10813_ _03750_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__clkbuf_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _07316_ _07317_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__nand2_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _04568_ _04569_ _04570_ _04225_ _04209_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__o221a_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16320_ _08282_ _07959_ vssd1 vssd1 vccd1 vccd1 _08965_ sky130_fd_sc_hd__nor2_1
X_19591__47 clknet_1_0__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__inv_2
XFILLER_186_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13532_ _06235_ _06268_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__xnor2_1
X_10744_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _03706_ vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16251_ _08895_ _08579_ vssd1 vssd1 vccd1 vccd1 _08896_ sky130_fd_sc_hd__or2_1
XFILLER_174_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13463_ _06160_ _06162_ _06163_ _06164_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__a22o_1
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10675_ rbzero.tex_g1\[19\] rbzero.tex_g1\[20\] _03669_ vssd1 vssd1 vccd1 vccd1 _03678_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15202_ _04028_ vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__buf_4
X_12414_ _05146_ _04325_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__nor2_1
XFILLER_185_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16182_ _08820_ _08826_ vssd1 vssd1 vccd1 vccd1 _08827_ sky130_fd_sc_hd__xor2_1
XFILLER_12_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13394_ _06129_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__xnor2_1
XFILLER_138_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15133_ _07786_ _07787_ _07783_ _07784_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__a211o_1
X_12345_ net42 _05103_ _05085_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__a31o_1
XFILLER_182_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15064_ _07720_ _07725_ _04033_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__mux2_1
X_19941_ _03231_ _03234_ _02714_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__o21a_1
X_12276_ net68 _05043_ _05044_ _04323_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__a22o_1
XFILLER_181_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14015_ _06744_ _06751_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__xnor2_1
X_11227_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__inv_2
X_19872_ rbzero.pov.ready_buffer\[71\] _03146_ _03180_ _03181_ _03155_ vssd1 vssd1
+ vccd1 vccd1 _03182_ sky130_fd_sc_hd__o221a_1
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18823_ _02502_ _01553_ rbzero.wall_tracer.trackDistY\[3\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00616_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_150_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ rbzero.wall_tracer.mapX\[7\] rbzero.wall_tracer.mapX\[6\] rbzero.wall_tracer.mapX\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__or3_1
XFILLER_95_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15966_ _08584_ _08610_ vssd1 vssd1 vccd1 vccd1 _08611_ sky130_fd_sc_hd__nor2_1
X_18754_ _02442_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__clkbuf_1
X_11089_ rbzero.tex_b0\[15\] rbzero.tex_b0\[14\] _03887_ vssd1 vssd1 vccd1 vccd1 _03895_
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17705_ _10125_ _10133_ _10135_ vssd1 vssd1 vccd1 vccd1 _10270_ sky130_fd_sc_hd__and3_1
XFILLER_64_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14917_ _07591_ _07617_ _07619_ _07620_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__o211a_1
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18685_ _02375_ _02380_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__xnor2_1
X_15897_ _08512_ _08538_ vssd1 vssd1 vccd1 vccd1 _08542_ sky130_fd_sc_hd__nor2_1
XFILLER_48_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17636_ _09096_ _09480_ _09484_ _09368_ vssd1 vssd1 vccd1 vccd1 _10201_ sky130_fd_sc_hd__o22a_1
X_14848_ _07394_ _07464_ _07468_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__a21o_2
XFILLER_24_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17567_ _10130_ _10131_ _10132_ vssd1 vssd1 vccd1 vccd1 _10133_ sky130_fd_sc_hd__nand3_1
XFILLER_17_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14779_ _07511_ _07447_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__nor2_1
X_20123__155 clknet_1_1__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__inv_2
XFILLER_205_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16518_ rbzero.wall_tracer.visualWallDist\[7\] _04015_ vssd1 vssd1 vccd1 vccd1 _09162_
+ sky130_fd_sc_hd__nand2_4
X_19306_ rbzero.spi_registers.new_other\[8\] rbzero.spi_registers.spi_buffer\[8\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__mux2_1
XFILLER_177_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ _10062_ _10063_ vssd1 vssd1 vccd1 vccd1 _10064_ sky130_fd_sc_hd__or2_1
XFILLER_143_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16449_ _07941_ _08035_ _08046_ _08075_ vssd1 vssd1 vccd1 vccd1 _09093_ sky130_fd_sc_hd__o22ai_1
X_19237_ rbzero.spi_registers.new_vshift\[5\] _02763_ vssd1 vssd1 vccd1 vccd1 _02770_
+ sky130_fd_sc_hd__or2_1
XFILLER_192_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19168_ rbzero.othery\[4\] _02710_ _02725_ _02722_ vssd1 vssd1 vccd1 vccd1 _00738_
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18119_ _01751_ _01736_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__and2b_1
XFILLER_191_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19099_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.spi_buffer\[4\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__mux2_1
XFILLER_133_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21130_ clknet_leaf_94_i_clk _00899_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21061_ net151 _00830_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20012_ _04892_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__inv_2
XFILLER_28_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ clknet_leaf_19_i_clk _00683_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_55_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20845_ clknet_leaf_48_i_clk _00614_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20776_ clknet_leaf_61_i_clk _00545_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20098__132 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__inv_2
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10460_ rbzero.tex_r0\[58\] rbzero.tex_r0\[57\] _03558_ vssd1 vssd1 vccd1 vccd1 _03565_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10391_ _03526_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ _04843_ _04845_ _04849_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__a31o_2
XFILLER_191_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21328_ net249 _01097_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12061_ _04832_ _04834_ net68 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__a21oi_2
X_21259_ clknet_leaf_88_i_clk _01028_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-7\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11012_ rbzero.tex_b0\[52\] rbzero.tex_b0\[51\] _03854_ vssd1 vssd1 vccd1 vccd1 _03855_
+ sky130_fd_sc_hd__mux2_1
XFILLER_132_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15820_ _08120_ _08146_ _08168_ vssd1 vssd1 vccd1 vccd1 _08465_ sky130_fd_sc_hd__and3_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _08393_ _08395_ vssd1 vssd1 vccd1 vccd1 _08396_ sky130_fd_sc_hd__xnor2_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _05684_ _05689_ _05694_ _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__o211ai_4
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14702_ _07375_ _07435_ _07436_ _07438_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__a31o_1
XFILLER_205_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18470_ _08275_ _09484_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__nor2_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _04686_ _04689_ _04209_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__mux2_1
X_15682_ _08297_ _08326_ vssd1 vssd1 vccd1 vccd1 _08327_ sky130_fd_sc_hd__xor2_4
XFILLER_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12894_ _05454_ _05630_ _05561_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__mux2_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17421_ _05210_ rbzero.wall_tracer.stepDistX\[9\] vssd1 vssd1 vccd1 vccd1 _09988_
+ sky130_fd_sc_hd__nand2_1
XFILLER_166_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _05893_ _07369_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__nand2_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _04266_ _04621_ _04229_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__o21a_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _09638_ _09652_ _09650_ vssd1 vssd1 vccd1 vccd1 _09919_ sky130_fd_sc_hd__a21o_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14564_ _07295_ _07300_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__and2b_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11776_ _04253_ _04549_ _04553_ _04119_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a211o_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16303_ _08945_ _08947_ vssd1 vssd1 vccd1 vccd1 _08948_ sky130_fd_sc_hd__xnor2_1
X_13515_ _06236_ _06250_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__or2_1
XFILLER_207_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10727_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _03624_ vssd1 vssd1 vccd1 vccd1 _03705_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17283_ _09846_ _09848_ _09847_ vssd1 vssd1 vccd1 vccd1 _09856_ sky130_fd_sc_hd__a21boi_1
X_14495_ _07220_ _07226_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__nor2_1
X_19022_ _02642_ vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16234_ _08877_ _08878_ vssd1 vssd1 vccd1 vccd1 _08879_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13446_ _06177_ _06178_ _06182_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10658_ _03646_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__clkbuf_4
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16165_ _08692_ _08718_ _08809_ vssd1 vssd1 vccd1 vccd1 _08810_ sky130_fd_sc_hd__a21oi_2
XFILLER_154_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13377_ _05995_ _06113_ _05846_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__a21o_1
X_10589_ _03632_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15116_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.debug_overlay.vplaneX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__and2_1
XFILLER_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12328_ _05087_ net66 _05095_ net30 vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__a211o_1
XFILLER_170_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16096_ _08733_ _08726_ vssd1 vssd1 vccd1 vccd1 _08741_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15047_ _04462_ rbzero.wall_tracer.rayAddendX\[-3\] vssd1 vssd1 vccd1 vccd1 _07710_
+ sky130_fd_sc_hd__nor2_1
X_19924_ rbzero.debug_overlay.playerY\[1\] _03216_ _03220_ vssd1 vssd1 vccd1 vccd1
+ _03221_ sky130_fd_sc_hd__a21o_1
X_12259_ _05021_ _04325_ vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__nor2_1
XFILLER_170_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19855_ _03145_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__nand2_1
XFILLER_69_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18806_ _02486_ _02487_ _02481_ _02483_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a211o_1
X_20398__23 clknet_1_0__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__inv_2
XFILLER_56_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19786_ rbzero.pov.spi_buffer\[66\] rbzero.pov.spi_buffer\[67\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03122_ sky130_fd_sc_hd__mux2_1
X_16998_ _09636_ _09637_ vssd1 vssd1 vccd1 vccd1 _09638_ sky130_fd_sc_hd__and2_1
XFILLER_96_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18737_ _02427_ vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15949_ _07990_ _08515_ vssd1 vssd1 vccd1 vccd1 _08594_ sky130_fd_sc_hd__nand2_2
XFILLER_184_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18668_ _02350_ _02363_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17619_ _09906_ _10183_ vssd1 vssd1 vccd1 vccd1 _10184_ sky130_fd_sc_hd__nor2_1
XFILLER_197_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18599_ _02179_ _02182_ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20630_ clknet_leaf_15_i_clk _00414_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20561_ rbzero.traced_texVinit\[4\] _03443_ _09771_ _03444_ vssd1 vssd1 vccd1 vccd1
+ _01412_ sky130_fd_sc_hd__a22o_1
XFILLER_165_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20492_ _03384_ _03388_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__nand2_1
XFILLER_164_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21113_ net203 _00882_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21044_ clknet_leaf_81_i_clk _00813_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11630_ _04244_ _04400_ _04408_ _04116_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__a31o_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20828_ clknet_leaf_50_i_clk _00597_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11561_ _04247_ _04334_ _04335_ _04339_ _04254_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__o221a_1
X_20759_ clknet_leaf_46_i_clk _00528_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_183_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13300_ _06030_ _06035_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__nand3b_1
X_10512_ _03592_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14280_ _06705_ _07016_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__xnor2_2
XFILLER_196_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11492_ _04271_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__buf_4
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13231_ _05929_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__or2_1
XFILLER_100_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10443_ _03475_ _03478_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__nand2_2
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13162_ _05834_ _05895_ _05898_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_opt_10_1_i_clk clknet_opt_10_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_10_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10374_ rbzero.tex_r1\[32\] rbzero.tex_r1\[33\] _03516_ vssd1 vssd1 vccd1 vccd1 _03518_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12113_ _04883_ _04884_ _04840_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__mux2_1
XFILLER_123_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17970_ _10294_ _10185_ _01550_ _01672_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a31oi_2
XFILLER_123_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13093_ _05733_ _05705_ _05792_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__mux2_1
X_20152__181 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__inv_2
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16921_ _09560_ _09561_ vssd1 vssd1 vccd1 vccd1 _09562_ sky130_fd_sc_hd__xor2_1
X_12044_ rbzero.row_render.wall\[0\] rbzero.row_render.wall\[1\] vssd1 vssd1 vccd1
+ vccd1 _04818_ sky130_fd_sc_hd__xnor2_2
XFILLER_105_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16852_ _09356_ _09357_ vssd1 vssd1 vccd1 vccd1 _09493_ sky130_fd_sc_hd__nand2_1
XFILLER_133_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15803_ _08446_ _08447_ vssd1 vssd1 vccd1 vccd1 _08448_ sky130_fd_sc_hd__xnor2_2
XFILLER_168_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16783_ _09423_ _09424_ vssd1 vssd1 vccd1 vccd1 _09425_ sky130_fd_sc_hd__nor2_1
X_19571_ clknet_1_0__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__buf_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13995_ _06731_ _06700_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__nor2_1
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18522_ _01922_ _02219_ _02112_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__o21a_1
X_15734_ _08303_ _08378_ vssd1 vssd1 vccd1 vccd1 _08379_ sky130_fd_sc_hd__xnor2_2
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12946_ _05674_ _05682_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__or2_2
XFILLER_206_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18453_ _02045_ _02150_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__nand2_1
X_15665_ _08308_ _08309_ vssd1 vssd1 vccd1 vccd1 _08310_ sky130_fd_sc_hd__xnor2_2
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _04030_ _05337_ _05344_ _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__a31o_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _09958_ _09970_ vssd1 vssd1 vccd1 vccd1 _09971_ sky130_fd_sc_hd__xnor2_1
X_14616_ _05931_ _07352_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__or2_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _02081_ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__and2_1
X_11828_ rbzero.tex_g1\[57\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__and3_1
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15596_ _08229_ _08240_ vssd1 vssd1 vccd1 vccd1 _08241_ sky130_fd_sc_hd__xor2_4
XFILLER_18_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _09889_ _09901_ _09902_ _09780_ vssd1 vssd1 vccd1 vccd1 _09903_ sky130_fd_sc_hd__a31o_1
X_14547_ _07279_ _07283_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__xnor2_1
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11759_ _04534_ _04535_ _04536_ _04224_ _04123_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__o221a_1
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17266_ _09838_ _09839_ _09840_ vssd1 vssd1 vccd1 vccd1 _09841_ sky130_fd_sc_hd__nor3_1
XFILLER_201_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14478_ _07213_ _07214_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__nor2_1
XFILLER_174_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16217_ _08854_ _08861_ vssd1 vssd1 vccd1 vccd1 _08862_ sky130_fd_sc_hd__xor2_1
XFILLER_128_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19005_ _02633_ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13429_ _06158_ _06165_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__xnor2_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17197_ _09777_ _09778_ _09779_ _09781_ rbzero.wall_tracer.mapX\[6\] vssd1 vssd1
+ vccd1 vccd1 _00571_ sky130_fd_sc_hd__a32o_1
X_20235__256 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__inv_2
X_16148_ _08284_ _08579_ _08727_ vssd1 vssd1 vccd1 vccd1 _08793_ sky130_fd_sc_hd__nor3_1
XFILLER_154_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079_ _08684_ _08686_ vssd1 vssd1 vccd1 vccd1 _08724_ sky130_fd_sc_hd__xnor2_1
X_19907_ _05190_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__buf_6
XFILLER_60_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19838_ rbzero.debug_overlay.playerX\[-5\] _03155_ vssd1 vssd1 vccd1 vccd1 _03156_
+ sky130_fd_sc_hd__or2_1
XFILLER_151_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput1 i_debug_vec_overlay vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_6
X_19769_ rbzero.pov.spi_buffer\[58\] rbzero.pov.spi_buffer\[59\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03113_ sky130_fd_sc_hd__mux2_1
XFILLER_65_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21662_ clknet_leaf_78_i_clk _01431_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20613_ _02721_ _03470_ _03471_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__and3_1
X_21593_ net134 _01362_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20544_ _09750_ _03433_ _03434_ _03250_ rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1
+ _01405_ sky130_fd_sc_hd__a32o_1
XFILLER_192_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20475_ rbzero.texV\[-2\] _03175_ _03332_ _03376_ vssd1 vssd1 vccd1 vccd1 _01394_
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21027_ clknet_leaf_4_i_clk _00796_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_other
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_142_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12800_ _05539_ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__or2b_1
X_13780_ _06514_ _06513_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__xnor2_1
X_10992_ _03844_ vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__and2_1
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20392__18 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__inv_2
XFILLER_128_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15450_ _05197_ _08094_ vssd1 vssd1 vccd1 vccd1 _08095_ sky130_fd_sc_hd__or2_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _03999_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__inv_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _07136_ _07137_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__xnor2_1
X_11613_ _04211_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__buf_6
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15381_ _08013_ _08025_ vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__or2b_1
X_12593_ _05289_ _05295_ _05303_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__nand3_1
XFILLER_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _04417_ _09748_ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__nor2_1
X_14332_ _06675_ _06708_ _07064_ _07068_ vssd1 vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__o31a_1
XFILLER_184_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11544_ _04314_ _04321_ _04323_ _04020_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__a211o_2
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ _09689_ _09690_ vssd1 vssd1 vccd1 vccd1 _09691_ sky130_fd_sc_hd__or2b_1
XFILLER_167_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14263_ _06698_ _06726_ _06672_ _06729_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__o31a_1
X_11475_ _04219_ _04249_ _04252_ _04254_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__o211a_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03289_ clknet_0__03289_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03289_
+ sky130_fd_sc_hd__clkbuf_16
X_16002_ _08644_ _08645_ _08646_ vssd1 vssd1 vccd1 vccd1 _08647_ sky130_fd_sc_hd__a21oi_1
X_13214_ _05826_ _05893_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10426_ rbzero.tex_r1\[7\] rbzero.tex_r1\[8\] _03538_ vssd1 vssd1 vccd1 vccd1 _03545_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14194_ _06924_ _06930_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__xnor2_1
XFILLER_136_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13145_ _05710_ _05640_ _05648_ _05687_ _05778_ _05792_ vssd1 vssd1 vccd1 vccd1 _05882_
+ sky130_fd_sc_hd__mux4_1
X_10357_ rbzero.tex_r1\[40\] rbzero.tex_r1\[41\] _03505_ vssd1 vssd1 vccd1 vccd1 _03509_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _01611_ _01655_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__xor2_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _05754_ _05797_ _05700_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a21oi_1
X_16904_ _07959_ _09126_ vssd1 vssd1 vccd1 vccd1 _09545_ sky130_fd_sc_hd__nor2_2
X_12027_ _04800_ _04801_ _04218_ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__mux2_1
X_17884_ _09391_ _09359_ _01463_ _10205_ _01462_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__o32a_1
XFILLER_66_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16835_ _09474_ _09475_ vssd1 vssd1 vccd1 vccd1 _09476_ sky130_fd_sc_hd__nor2_1
XFILLER_20_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19554_ _03022_ _03023_ _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__and3b_1
XFILLER_20_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16766_ _09278_ _09280_ _09281_ _09277_ vssd1 vssd1 vccd1 vccd1 _09408_ sky130_fd_sc_hd__a22oi_2
X_13978_ _06714_ _06674_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18505_ _02200_ _02201_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__and2_1
XFILLER_94_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15717_ _07967_ _08097_ vssd1 vssd1 vccd1 vccd1 _08362_ sky130_fd_sc_hd__or2_1
X_12929_ _05650_ _05655_ _05664_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16697_ rbzero.wall_tracer.texu\[2\] _09085_ vssd1 vssd1 vccd1 vccd1 _09340_ sky130_fd_sc_hd__or2_1
X_19485_ _02963_ _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nand2_1
XFILLER_94_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18436_ _02132_ _02133_ _02134_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__o21ai_1
XFILLER_181_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15648_ _07996_ _07958_ vssd1 vssd1 vccd1 vccd1 _08293_ sky130_fd_sc_hd__nor2_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18367_ _01474_ _09350_ _01934_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__nor3_1
X_15579_ _07970_ _08222_ _08223_ _07951_ vssd1 vssd1 vccd1 vccd1 _08224_ sky130_fd_sc_hd__a31o_2
XFILLER_159_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17318_ _09887_ vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__clkbuf_1
X_18298_ _01977_ _01997_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__xnor2_2
XFILLER_174_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17249_ _08944_ _08948_ _04016_ vssd1 vssd1 vccd1 vccd1 _09826_ sky130_fd_sc_hd__o21ai_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20260_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__buf_1
XFILLER_190_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21645_ clknet_leaf_29_i_clk _01414_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21576_ net497 _01345_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[27\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_50 _09859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_72 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_83 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20527_ rbzero.texV\[6\] _03327_ _03332_ _03420_ vssd1 vssd1 vccd1 vccd1 _01402_
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20218__240 clknet_1_0__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__inv_2
XFILLER_119_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11260_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__inv_2
X_20458_ rbzero.traced_texa\[-4\] rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1 _03362_
+ sky130_fd_sc_hd__nor2_1
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11191_ rbzero.map_rom.f4 rbzero.map_rom.f3 _03973_ _03979_ vssd1 vssd1 vccd1 vccd1
+ _03980_ sky130_fd_sc_hd__a31o_1
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14950_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.trackDistX\[8\] _05278_
+ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__mux2_1
XFILLER_87_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13901_ _06619_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__xnor2_2
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14881_ _03969_ _04017_ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__nor2_2
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16620_ _09241_ _09242_ _09262_ vssd1 vssd1 vccd1 vccd1 _09263_ sky130_fd_sc_hd__a21o_1
X_13832_ _05974_ _06161_ _05940_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__or3_1
XFILLER_78_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20264__282 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__inv_2
XFILLER_28_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16551_ rbzero.debug_overlay.playerY\[-5\] _07895_ vssd1 vssd1 vccd1 vccd1 _09195_
+ sky130_fd_sc_hd__or2_1
X_13763_ _06491_ _06492_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__and2_1
X_10975_ _03835_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _07945_ vssd1 vssd1 vccd1 vccd1 _08147_ sky130_fd_sc_hd__buf_4
X_12714_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__nand2_1
XFILLER_44_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16482_ _08189_ vssd1 vssd1 vccd1 vccd1 _09126_ sky130_fd_sc_hd__clkbuf_4
X_19270_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_floor\[5\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__mux2_1
X_13694_ _06429_ _06430_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__xor2_1
XFILLER_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18221_ _01920_ _01825_ _01823_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15433_ rbzero.debug_overlay.playerX\[-2\] vssd1 vssd1 vccd1 vccd1 _08078_ sky130_fd_sc_hd__inv_2
XFILLER_176_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12645_ _05396_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18152_ _01838_ _01852_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15364_ _08008_ _07932_ vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__nor2_1
XFILLER_8_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12576_ _05324_ _05325_ _05328_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__nand3_1
XFILLER_15_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17103_ _09599_ vssd1 vssd1 vccd1 vccd1 _09743_ sky130_fd_sc_hd__inv_2
X_14315_ _06997_ _06726_ _07051_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__o21a_1
X_18083_ _01686_ _01784_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__xor2_1
X_11527_ _04247_ _04302_ _04303_ _04305_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__o221a_1
XFILLER_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15295_ _07938_ _07939_ vssd1 vssd1 vccd1 vccd1 _07940_ sky130_fd_sc_hd__or2_1
XFILLER_117_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17034_ _09103_ vssd1 vssd1 vccd1 vccd1 _09674_ sky130_fd_sc_hd__clkbuf_4
XFILLER_176_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14246_ _06944_ _06969_ _06975_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__and3_1
X_11458_ rbzero.tex_r0\[55\] _04221_ _04222_ _04219_ vssd1 vssd1 vccd1 vccd1 _04238_
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10409_ rbzero.tex_r1\[15\] rbzero.tex_r1\[16\] _03527_ vssd1 vssd1 vccd1 vccd1 _03536_
+ sky130_fd_sc_hd__mux2_1
X_14177_ _06905_ _06913_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__nand2_1
X_11389_ _04161_ _04022_ gpout0.hpos\[3\] _04162_ _04168_ vssd1 vssd1 vccd1 vccd1
+ _04169_ sky130_fd_sc_hd__a221o_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _05798_ _05864_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__nor2_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ rbzero.pov.spi_buffer\[25\] rbzero.pov.ready_buffer\[25\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02623_ sky130_fd_sc_hd__mux2_1
XFILLER_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _01636_ _01637_ _01638_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__nand3_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _05775_ _05788_ _05789_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__nor3_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20347__357 clknet_1_0__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__inv_2
XFILLER_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17867_ _01561_ _01562_ _01568_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__and3_1
XFILLER_39_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16818_ _09459_ _08067_ _07895_ vssd1 vssd1 vccd1 vccd1 _09460_ sky130_fd_sc_hd__mux2_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17798_ _01500_ _01501_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__xnor2_2
XFILLER_207_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19537_ rbzero.wall_tracer.rayAddendY\[10\] _07695_ _07830_ _03012_ vssd1 vssd1 vccd1
+ vccd1 _03013_ sky130_fd_sc_hd__o2bb2a_1
X_16749_ _09245_ vssd1 vssd1 vccd1 vccd1 _09391_ sky130_fd_sc_hd__clkbuf_4
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03037_ clknet_0__03037_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03037_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19468_ _02904_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02949_
+ sky130_fd_sc_hd__or2_1
XFILLER_179_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18419_ _02116_ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19399_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.debug_overlay.vplaneY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__nor2_1
X_21430_ net351 _01199_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21361_ net282 _01130_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20092__127 clknet_1_0__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__inv_2
XFILLER_174_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21292_ clknet_leaf_3_i_clk _01061_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_72_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_87_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10760_ rbzero.tex_g0\[44\] rbzero.tex_g0\[43\] _03718_ vssd1 vssd1 vccd1 vccd1 _03723_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10691_ _03686_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_10_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_139_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12430_ net71 rbzero.wall_tracer.state\[7\] _05190_ vssd1 vssd1 vccd1 vccd1 _05192_
+ sky130_fd_sc_hd__and3_1
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21628_ clknet_leaf_46_i_clk _01397_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12361_ _05101_ _05126_ _05128_ _05085_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_139_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21559_ net480 _01328_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14100_ _06822_ _06835_ _06836_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__a21boi_1
XFILLER_10_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11312_ _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__inv_2
X_15080_ _07728_ _07734_ _07740_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__a21o_1
XFILLER_10_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12292_ net25 _05052_ _05060_ _05034_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__o211a_1
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14031_ _06766_ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__nand2_1
X_11243_ rbzero.wall_tracer.state\[14\] _04021_ _04026_ vssd1 vssd1 vccd1 vccd1 _04027_
+ sky130_fd_sc_hd__and3_2
XFILLER_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11174_ rbzero.otherx\[3\] _03936_ _03919_ rbzero.otherx\[0\] vssd1 vssd1 vccd1 vccd1
+ _03963_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_122_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18770_ _02456_ vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15982_ _08626_ _08039_ _08040_ vssd1 vssd1 vccd1 vccd1 _08627_ sky130_fd_sc_hd__and3_1
XFILLER_94_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17721_ _10156_ _10158_ vssd1 vssd1 vccd1 vccd1 _10286_ sky130_fd_sc_hd__nor2_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14933_ _07621_ _07630_ _07631_ _07620_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__o211a_1
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17652_ _08445_ _08418_ vssd1 vssd1 vccd1 vccd1 _10217_ sky130_fd_sc_hd__nand2_1
X_14864_ _07580_ vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16603_ _07932_ _08129_ _08047_ _09245_ vssd1 vssd1 vccd1 vccd1 _09246_ sky130_fd_sc_hd__o22ai_1
XFILLER_91_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13815_ _06548_ _06549_ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__o21ai_1
X_17583_ _09994_ _10002_ vssd1 vssd1 vccd1 vccd1 _10149_ sky130_fd_sc_hd__or2_1
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14795_ _07473_ _07478_ vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__nand2_1
XFILLER_17_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19322_ _02817_ vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__clkbuf_1
X_16534_ _09161_ _09166_ _09177_ vssd1 vssd1 vccd1 vccd1 _09178_ sky130_fd_sc_hd__or3b_1
XFILLER_32_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13746_ _06469_ _06471_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__nand2_1
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10958_ _03826_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19253_ _02779_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__clkbuf_1
X_16465_ _09098_ _09108_ vssd1 vssd1 vccd1 vccd1 _09109_ sky130_fd_sc_hd__xnor2_1
X_13677_ _06398_ _06412_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__nor2_1
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10889_ _03790_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__clkbuf_1
X_18204_ _01903_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__or2_1
X_12628_ rbzero.map_rom.b6 _05374_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__and2_1
X_15416_ _07933_ _08060_ _07903_ vssd1 vssd1 vccd1 vccd1 _08061_ sky130_fd_sc_hd__a21o_1
X_16396_ _08161_ _08431_ vssd1 vssd1 vccd1 vccd1 _09041_ sky130_fd_sc_hd__nor2_1
X_19184_ rbzero.spi_registers.new_leak\[3\] _02733_ vssd1 vssd1 vccd1 vccd1 _02737_
+ sky130_fd_sc_hd__or2_1
XFILLER_185_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18135_ _01826_ _01835_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__nand2_1
X_15347_ _07545_ _07991_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _07992_
+ sky130_fd_sc_hd__mux2_2
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12559_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__nor2_1
XFILLER_184_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18066_ _01754_ _01647_ _01766_ _01767_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__a211o_1
XFILLER_145_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15278_ _07922_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__clkbuf_2
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17017_ _09617_ _09656_ vssd1 vssd1 vccd1 vccd1 _09657_ sky130_fd_sc_hd__xnor2_2
X_14229_ _06964_ _06965_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__and2_1
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ rbzero.pov.spi_buffer\[17\] rbzero.pov.ready_buffer\[17\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02614_ sky130_fd_sc_hd__mux2_1
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17919_ _01619_ _01621_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__and2_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18899_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\] _02560_
+ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__and3_1
XFILLER_78_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20930_ clknet_leaf_26_i_clk _00699_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20861_ clknet_leaf_0_i_clk _00630_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20792_ clknet_leaf_28_i_clk _00561_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20100__134 clknet_1_1__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__inv_2
XFILLER_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21413_ net334 _01182_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_185_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21344_ net265 _01113_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21275_ clknet_leaf_93_i_clk _01044_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ rbzero.tex_b0\[59\] rbzero.tex_b0\[58\] _04263_ vssd1 vssd1 vccd1 vccd1 _04706_
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11861_ rbzero.tex_g1\[7\] rbzero.tex_g1\[6\] _04336_ vssd1 vssd1 vccd1 vccd1 _04638_
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _06293_ _06296_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__xnor2_1
XFILLER_14_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10812_ rbzero.tex_g0\[19\] rbzero.tex_g0\[18\] _03740_ vssd1 vssd1 vccd1 vccd1 _03750_
+ sky130_fd_sc_hd__mux2_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _07273_ _07278_ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__xor2_2
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _04262_ vssd1 vssd1 vccd1 vccd1 _04570_
+ sky130_fd_sc_hd__mux2_1
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _06253_ _06267_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__xnor2_1
XFILLER_159_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10743_ _03713_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16250_ _08283_ vssd1 vssd1 vccd1 vccd1 _08895_ sky130_fd_sc_hd__clkbuf_4
XFILLER_51_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _05752_ _06153_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__nand2_1
X_10674_ _03677_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20376__383 clknet_1_0__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__inv_2
XFILLER_185_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15201_ _07851_ _07852_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__or2_1
XFILLER_40_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12413_ _05146_ net61 _05179_ net36 vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__o211a_1
X_16181_ _08816_ _08821_ _08825_ _08822_ vssd1 vssd1 vccd1 vccd1 _08826_ sky130_fd_sc_hd__o31a_1
XFILLER_199_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13393_ _06039_ _06048_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20075__111 clknet_1_0__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__inv_2
X_15132_ _07788_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__inv_2
X_12344_ _05082_ _05083_ _04021_ _05085_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__and4_1
XFILLER_166_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15063_ _07723_ _07724_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__xnor2_1
X_19940_ rbzero.pov.ready_buffer\[57\] _03164_ _03233_ vssd1 vssd1 vccd1 vccd1 _03234_
+ sky130_fd_sc_hd__o21a_1
X_12275_ net21 net20 vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__nor2_2
XFILLER_141_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14014_ _06745_ _06750_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__xnor2_2
X_11226_ _04011_ _04007_ _03478_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__a21bo_1
XFILLER_107_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19871_ rbzero.debug_overlay.playerX\[3\] _03176_ _02822_ vssd1 vssd1 vccd1 vccd1
+ _03181_ sky130_fd_sc_hd__a21o_1
XFILLER_96_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18822_ _09889_ _02501_ _02399_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a21boi_1
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11157_ _03940_ _03941_ _03943_ _03944_ _03945_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a221o_1
XFILLER_110_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18753_ rbzero.wall_tracer.trackDistY\[-6\] _02440_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02442_ sky130_fd_sc_hd__mux2_1
X_15965_ _08492_ _08566_ _08583_ vssd1 vssd1 vccd1 vccd1 _08610_ sky130_fd_sc_hd__and3_1
XFILLER_49_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11088_ _03894_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__clkbuf_1
X_17704_ _10265_ _10268_ vssd1 vssd1 vccd1 vccd1 _10269_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14916_ _04035_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__buf_2
X_18684_ _02377_ _02379_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__xnor2_1
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15896_ _08509_ _08540_ vssd1 vssd1 vccd1 vccd1 _08541_ sky130_fd_sc_hd__nor2_1
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17635_ _09096_ _09480_ _09484_ vssd1 vssd1 vccd1 vccd1 _10200_ sky130_fd_sc_hd__or3_1
XFILLER_1_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14847_ _07567_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17566_ _09117_ _10129_ vssd1 vssd1 vccd1 vccd1 _10132_ sky130_fd_sc_hd__nor2_1
XFILLER_189_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14778_ _07486_ _07433_ vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__nand2_1
XFILLER_95_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19305_ _02808_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__clkbuf_1
X_16517_ rbzero.wall_tracer.visualWallDist\[7\] _04015_ _09030_ _08416_ vssd1 vssd1
+ vccd1 vccd1 _09161_ sky130_fd_sc_hd__and4_1
XFILLER_17_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1055 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13729_ _06453_ _06452_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__or2b_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17497_ _09368_ _09217_ _09929_ _09927_ vssd1 vssd1 vccd1 vccd1 _10063_ sky130_fd_sc_hd__o31a_1
XFILLER_108_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19236_ rbzero.spi_registers.vshift\[4\] _02762_ _02769_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00762_ sky130_fd_sc_hd__o211a_1
XFILLER_177_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16448_ _07941_ _08075_ _08035_ _08046_ vssd1 vssd1 vccd1 vccd1 _09092_ sky130_fd_sc_hd__or4_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19167_ rbzero.spi_registers.new_other\[4\] _02712_ vssd1 vssd1 vccd1 vccd1 _02725_
+ sky130_fd_sc_hd__or2_1
XFILLER_173_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16379_ _08327_ _08370_ _09023_ vssd1 vssd1 vccd1 vccd1 _09024_ sky130_fd_sc_hd__a21oi_4
XFILLER_157_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18118_ _01715_ _01730_ _01818_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__a21o_1
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19098_ _02682_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__clkbuf_1
XFILLER_172_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18049_ _01743_ _01750_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__xnor2_1
XFILLER_28_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21060_ net150 _00829_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20011_ _04892_ _04992_ _04884_ _04883_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__or4bb_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20913_ clknet_leaf_19_i_clk _00682_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20844_ clknet_leaf_61_i_clk _00613_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20775_ clknet_leaf_39_i_clk _00544_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10390_ rbzero.tex_r1\[24\] rbzero.tex_r1\[25\] _03516_ vssd1 vssd1 vccd1 vccd1 _03526_
+ sky130_fd_sc_hd__mux2_1
XFILLER_135_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21327_ net248 _01096_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12060_ _03474_ _04820_ _04833_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__a21o_1
XFILLER_172_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21258_ clknet_leaf_90_i_clk _01027_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_145_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11011_ _03717_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__clkbuf_4
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21189_ clknet_leaf_23_i_clk _00958_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _08394_ _08315_ vssd1 vssd1 vccd1 vccd1 _08395_ sky130_fd_sc_hd__xor2_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12962_ _05695_ _05673_ _05696_ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__or4_2
XFILLER_86_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14701_ _05963_ _07437_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__and2_1
X_11913_ _04687_ _04688_ _04139_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__mux2_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15681_ _08313_ _08324_ _08325_ vssd1 vssd1 vccd1 vccd1 _08326_ sky130_fd_sc_hd__a21oi_2
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12893_ _04031_ _05329_ _05330_ _05629_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__a31o_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _09117_ _09693_ vssd1 vssd1 vccd1 vccd1 _09987_ sky130_fd_sc_hd__nor2_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ rbzero.tex_g1\[35\] rbzero.tex_g1\[34\] _04350_ vssd1 vssd1 vccd1 vccd1 _04621_
+ sky130_fd_sc_hd__mux2_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14632_ _07367_ _07315_ _07368_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17351_ _09908_ _09917_ vssd1 vssd1 vccd1 vccd1 _09918_ sky130_fd_sc_hd__xor2_4
X_14563_ _07297_ _07299_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__nor2_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _04224_ _04550_ _04551_ _04552_ _04141_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__o221a_1
XFILLER_53_1206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _08941_ _08811_ _08946_ vssd1 vssd1 vccd1 vccd1 _08947_ sky130_fd_sc_hd__a21oi_1
XFILLER_202_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10726_ _03704_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13514_ _06236_ _06250_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__nand2_1
XFILLER_147_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14494_ _07229_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__and2b_1
X_17282_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _09855_ sky130_fd_sc_hd__and2_1
XFILLER_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19021_ rbzero.pov.spi_buffer\[42\] rbzero.pov.ready_buffer\[42\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02642_ sky130_fd_sc_hd__mux2_1
X_16233_ _08830_ _08868_ vssd1 vssd1 vccd1 vccd1 _08878_ sky130_fd_sc_hd__xnor2_1
X_13445_ _06179_ _06181_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__xnor2_1
X_10657_ _03668_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13376_ _05889_ _05900_ _05910_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__a21o_1
X_16164_ _08693_ _08717_ vssd1 vssd1 vccd1 vccd1 _08809_ sky130_fd_sc_hd__nor2_1
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10588_ rbzero.tex_g1\[60\] rbzero.tex_g1\[61\] _03549_ vssd1 vssd1 vccd1 vccd1 _03632_
+ sky130_fd_sc_hd__mux2_1
X_12327_ _05087_ _04325_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__nor2_1
XFILLER_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15115_ _07758_ _07761_ _07771_ _03912_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__a31o_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16095_ _08697_ _08712_ vssd1 vssd1 vccd1 vccd1 _08740_ sky130_fd_sc_hd__xnor2_1
XFILLER_108_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15046_ rbzero.debug_overlay.vplaneX\[-7\] _07705_ vssd1 vssd1 vccd1 vccd1 _07709_
+ sky130_fd_sc_hd__nand2_1
X_19923_ rbzero.debug_overlay.playerY\[1\] _03216_ _03145_ vssd1 vssd1 vccd1 vccd1
+ _03220_ sky130_fd_sc_hd__o21ai_1
X_12258_ net25 vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__inv_2
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11209_ rbzero.wall_tracer.state\[1\] _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__nand2_1
X_19854_ rbzero.debug_overlay.playerX\[0\] _08028_ vssd1 vssd1 vccd1 vccd1 _03167_
+ sky130_fd_sc_hd__or2_1
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18805_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__nand2_1
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19785_ _03121_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16997_ _09626_ _09635_ vssd1 vssd1 vccd1 vccd1 _09637_ sky130_fd_sc_hd__or2_1
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18736_ rbzero.wall_tracer.trackDistY\[-8\] _02426_ _02399_ vssd1 vssd1 vccd1 vccd1
+ _02427_ sky130_fd_sc_hd__mux2_1
XFILLER_83_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15948_ _08591_ _08592_ vssd1 vssd1 vccd1 vccd1 _08593_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18667_ _02351_ _02362_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__xnor2_1
XFILLER_149_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15879_ _08520_ _08521_ vssd1 vssd1 vccd1 vccd1 _08524_ sky130_fd_sc_hd__and2_1
XFILLER_24_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17618_ _10165_ _10166_ _10026_ vssd1 vssd1 vccd1 vccd1 _10183_ sky130_fd_sc_hd__nand3b_1
XFILLER_184_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18598_ _02167_ _02168_ _02294_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a21boi_1
XFILLER_196_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17549_ _08283_ _09555_ vssd1 vssd1 vccd1 vccd1 _10115_ sky130_fd_sc_hd__nor2_1
XFILLER_189_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20560_ _09331_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__inv_2
XFILLER_20_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19219_ _09753_ _02758_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__and2_1
XFILLER_192_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20491_ rbzero.traced_texa\[1\] rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 _03390_
+ sky130_fd_sc_hd__nand2_1
XFILLER_30_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21112_ net202 _00881_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[52\] sky130_fd_sc_hd__dfxtp_1
X_20212__235 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__inv_2
XFILLER_87_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19618__71 clknet_1_0__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__inv_2
X_21043_ clknet_leaf_75_i_clk _00812_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_99_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19633__85 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__inv_2
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20827_ clknet_leaf_44_i_clk _00596_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11560_ rbzero.tex_r1\[10\] _04338_ _04304_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__a21o_1
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20758_ clknet_leaf_29_i_clk _00527_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.side
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10511_ rbzero.tex_r0\[34\] rbzero.tex_r0\[33\] _03591_ vssd1 vssd1 vccd1 vccd1 _03592_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ _04129_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__buf_6
XFILLER_137_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20689_ clknet_leaf_55_i_clk _00473_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13230_ _05826_ _05934_ _05965_ _05966_ _05928_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__o221a_1
XFILLER_108_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ _03553_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13161_ _05800_ _05896_ _05897_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__o21a_1
XFILLER_164_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10373_ _03517_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12112_ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__buf_2
XFILLER_3_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13092_ _05757_ _05773_ _05792_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__mux2_1
XFILLER_151_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12043_ _04811_ _04813_ _04815_ _04816_ _04005_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__a311o_1
X_16920_ _07598_ _09283_ _05210_ _09433_ vssd1 vssd1 vccd1 vccd1 _09561_ sky130_fd_sc_hd__or4_1
XFILLER_77_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20187__212 clknet_1_0__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__inv_2
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16851_ _09488_ _09491_ vssd1 vssd1 vccd1 vccd1 _09492_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15802_ _07974_ _08376_ vssd1 vssd1 vccd1 vccd1 _08447_ sky130_fd_sc_hd__or2_1
X_19570_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__buf_1
XFILLER_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16782_ _09418_ _09422_ vssd1 vssd1 vccd1 vccd1 _09424_ sky130_fd_sc_hd__nor2_1
XFILLER_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13994_ _06729_ _06730_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__nand2_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18521_ _02114_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__inv_2
XFILLER_206_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ _08275_ _08377_ vssd1 vssd1 vccd1 vccd1 _08378_ sky130_fd_sc_hd__nor2_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _05677_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__or2_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _08802_ _09668_ _01524_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a21oi_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15664_ _08282_ _08194_ vssd1 vssd1 vccd1 vccd1 _08309_ sky130_fd_sc_hd__nor2_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12876_ rbzero.wall_tracer.visualWallDist\[-3\] _05571_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05613_ sky130_fd_sc_hd__a21o_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _09963_ _09969_ vssd1 vssd1 vccd1 vccd1 _09970_ sky130_fd_sc_hd__xor2_2
XFILLER_178_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14615_ _07107_ _07349_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__a21o_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _02070_ _02080_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__or2_1
X_11827_ _04602_ _04603_ _04304_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__mux2_1
XFILLER_159_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _08237_ _08239_ vssd1 vssd1 vccd1 vccd1 _08240_ sky130_fd_sc_hd__nor2_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _09900_ _09893_ _09898_ _09899_ vssd1 vssd1 vccd1 vccd1 _09902_ sky130_fd_sc_hd__a211o_1
XFILLER_186_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11758_ rbzero.tex_g0\[1\] rbzero.tex_g0\[0\] _04341_ vssd1 vssd1 vccd1 vccd1 _04536_
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14546_ _07281_ _07282_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__nor2_1
XFILLER_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ rbzero.tex_g1\[3\] rbzero.tex_g1\[4\] _03691_ vssd1 vssd1 vccd1 vccd1 _03696_
+ sky130_fd_sc_hd__mux2_1
XFILLER_179_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17265_ _09830_ _09832_ _09831_ vssd1 vssd1 vccd1 vccd1 _09840_ sky130_fd_sc_hd__a21boi_1
XFILLER_197_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11689_ _04462_ _04463_ _04464_ rbzero.debug_overlay.vplaneX\[-4\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__a221o_1
X_14477_ _07211_ _07212_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__and2_1
X_19004_ rbzero.pov.spi_buffer\[34\] rbzero.pov.ready_buffer\[34\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02633_ sky130_fd_sc_hd__mux2_1
X_16216_ _08377_ _08062_ vssd1 vssd1 vccd1 vccd1 _08861_ sky130_fd_sc_hd__nor2_1
X_13428_ _06163_ _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17196_ _09780_ vssd1 vssd1 vccd1 vccd1 _09781_ sky130_fd_sc_hd__buf_6
X_16147_ _08787_ _08790_ _08791_ vssd1 vssd1 vccd1 vccd1 _08792_ sky130_fd_sc_hd__a21bo_1
X_13359_ _05941_ _05980_ _05990_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16078_ _08675_ _08720_ _08721_ _08722_ vssd1 vssd1 vccd1 vccd1 _08723_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_170_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15029_ _07682_ _07693_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__xnor2_1
X_19906_ rbzero.pov.ready_buffer\[49\] _02823_ _03192_ _03207_ vssd1 vssd1 vccd1 vccd1
+ _03208_ sky130_fd_sc_hd__a211o_1
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19837_ net38 _03137_ _02708_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__o21a_2
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 i_gpout0_sel[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_8
X_19768_ _03112_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18719_ _09863_ _02410_ _02411_ _09827_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__o31ai_1
X_19699_ _03076_ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03299_ _03299_ vssd1 vssd1 vccd1 vccd1 clknet_0__03299_ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21661_ clknet_leaf_76_i_clk _01430_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
X_20612_ gpout4.clk_div\[1\] gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__or2_1
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21592_ net133 _01361_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[43\] sky130_fd_sc_hd__dfxtp_1
X_20543_ _03430_ _03431_ _03432_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__nand3_1
XFILLER_138_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20474_ _03374_ _03375_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__xor2_1
XFILLER_192_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21026_ clknet_leaf_4_i_clk _00795_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10991_ rbzero.tex_b0\[62\] rbzero.tex_b0\[61\] _03843_ vssd1 vssd1 vccd1 vccd1 _03844_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ rbzero.wall_tracer.rayAddendX\[-4\] rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.rayAddendX\[-2\]
+ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__or4_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ rbzero.debug_overlay.playerX\[0\] _03919_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05410_ sky130_fd_sc_hd__mux2_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11612_ _04230_ _04386_ _04390_ _04242_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__a211o_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _06696_ _06708_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__nor2_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15380_ _08014_ _08023_ _08024_ vssd1 vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__a21bo_1
X_12592_ _05306_ _05343_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__xor2_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11543_ gpout0.vpos\[5\] _04322_ gpout0.vpos\[9\] vssd1 vssd1 vccd1 vccd1 _04323_
+ sky130_fd_sc_hd__a21o_4
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14331_ _06689_ _06663_ _07011_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__or3_1
XFILLER_195_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17050_ _09683_ _09688_ vssd1 vssd1 vccd1 vccd1 _09690_ sky130_fd_sc_hd__or2_1
X_14262_ _06996_ _06998_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__xnor2_1
X_11474_ _04253_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__buf_4
XFILLER_13_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13213_ _05848_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__inv_2
XFILLER_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16001_ _08642_ _08643_ vssd1 vssd1 vccd1 vccd1 _08646_ sky130_fd_sc_hd__and2b_1
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ _03544_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__clkbuf_1
X_14193_ _06895_ _06925_ _06929_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__a21bo_1
XFILLER_164_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ _05844_ _05880_ _05798_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__a21oi_2
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10356_ _03508_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17952_ _01653_ _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__xor2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13075_ _05802_ _05808_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__mux2_1
XFILLER_183_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16903_ _09409_ _09543_ vssd1 vssd1 vccd1 vccd1 _09544_ sky130_fd_sc_hd__xnor2_1
X_12026_ rbzero.tex_b1\[37\] rbzero.tex_b1\[36\] _04250_ vssd1 vssd1 vccd1 vccd1 _04801_
+ sky130_fd_sc_hd__mux2_1
X_17883_ _01584_ _01585_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__xor2_1
XFILLER_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16834_ _09379_ _09471_ _09473_ vssd1 vssd1 vccd1 vccd1 _09475_ sky130_fd_sc_hd__and3_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19553_ _03019_ _03025_ _03020_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__a21boi_1
XFILLER_20_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19612__66 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__inv_2
X_16765_ _09119_ _09270_ _09406_ vssd1 vssd1 vccd1 vccd1 _09407_ sky130_fd_sc_hd__a21bo_1
XFILLER_150_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13977_ _06240_ _06662_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__or2_1
XFILLER_59_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18504_ _02200_ _02201_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__nor2_1
XFILLER_111_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15716_ _08359_ _08360_ vssd1 vssd1 vccd1 vccd1 _08361_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19484_ _02905_ _04471_ rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1
+ _02964_ sky130_fd_sc_hd__or3b_1
X_12928_ _05650_ _05655_ _05664_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__or3_1
X_16696_ _09082_ _09338_ vssd1 vssd1 vccd1 vccd1 _09339_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18435_ _02017_ _02019_ _02018_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a21boi_1
XFILLER_62_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20241__261 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__inv_2
X_15647_ _08290_ _08291_ vssd1 vssd1 vccd1 vccd1 _08292_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _05477_ _05595_ _05560_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__mux2_4
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18366_ _02063_ _02064_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__nand2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15578_ _07893_ _05372_ vssd1 vssd1 vccd1 vccd1 _08223_ sky130_fd_sc_hd__or2_2
X_17317_ rbzero.wall_tracer.trackDistX\[-3\] _09886_ _05413_ vssd1 vssd1 vccd1 vccd1
+ _09887_ sky130_fd_sc_hd__mux2_1
X_14529_ _07264_ _07265_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__and2b_1
X_18297_ _01979_ _01996_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20159__188 clknet_1_1__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__inv_2
X_17248_ _09823_ _09821_ _09822_ _05531_ vssd1 vssd1 vccd1 vccd1 _09825_ sky130_fd_sc_hd__a31o_1
XFILLER_128_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17179_ rbzero.traced_texa\[7\] _09770_ _09769_ rbzero.wall_tracer.visualWallDist\[7\]
+ vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__a22o_1
XFILLER_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20324__336 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__inv_2
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_opt_10_0_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_10_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21644_ clknet_leaf_30_i_clk _01413_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_40 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21575_ net496 _01344_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_51 _10297_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_73 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20526_ _03418_ _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_84 net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20457_ _03272_ _03360_ _03361_ _03327_ rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1
+ _01391_ sky130_fd_sc_hd__a32o_1
X_20370__378 clknet_1_0__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__inv_2
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ _03919_ _03925_ _03976_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__a31o_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13900_ _06635_ _06636_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__xnor2_2
X_21009_ clknet_leaf_9_i_clk _00778_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_floor
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14880_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.trackDistX\[-12\]
+ _07592_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_i_clk clknet_1_1_1_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13831_ _06253_ _06267_ _06251_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__a21bo_1
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16550_ _09088_ _09193_ vssd1 vssd1 vccd1 vccd1 _09194_ sky130_fd_sc_hd__xnor2_4
X_20299__313 clknet_1_1__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__inv_2
X_10974_ rbzero.tex_b1\[5\] rbzero.tex_b1\[6\] _03828_ vssd1 vssd1 vccd1 vccd1 _03835_
+ sky130_fd_sc_hd__mux2_1
X_13762_ _06461_ _06458_ _06460_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__and3_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15501_ _08122_ _08145_ vssd1 vssd1 vccd1 vccd1 _08146_ sky130_fd_sc_hd__or2b_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12713_ _05442_ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__and2_1
XFILLER_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16481_ _09116_ _09124_ vssd1 vssd1 vccd1 vccd1 _09125_ sky130_fd_sc_hd__xnor2_2
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13693_ _05945_ _06409_ _06078_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__a21oi_1
X_18220_ _01822_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__inv_2
XFILLER_102_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15432_ rbzero.debug_overlay.playerX\[-2\] _08027_ vssd1 vssd1 vccd1 vccd1 _08077_
+ sky130_fd_sc_hd__xnor2_1
X_12644_ _05395_ rbzero.map_rom.a6 _05284_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__mux2_1
XFILLER_203_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18151_ _01850_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__nor2_1
XFILLER_197_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _05324_ _05325_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__a21o_1
X_15363_ _07945_ _08001_ _08006_ _08007_ vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__a22o_4
XFILLER_15_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17102_ _09739_ _09741_ vssd1 vssd1 vccd1 vccd1 _09742_ sky130_fd_sc_hd__xnor2_1
X_14314_ _06996_ _06998_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__nand2_1
XFILLER_89_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18082_ _01781_ _01783_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__xnor2_1
X_11526_ _04209_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__buf_4
XFILLER_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15294_ _05197_ rbzero.wall_tracer.stepDistX\[-5\] vssd1 vssd1 vccd1 vccd1 _07939_
+ sky130_fd_sc_hd__nor2_2
XFILLER_144_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17033_ _09669_ _09672_ vssd1 vssd1 vccd1 vccd1 _09673_ sky130_fd_sc_hd__xnor2_2
X_11457_ rbzero.tex_r0\[54\] _04214_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__and2_1
X_14245_ _06962_ _06979_ _06981_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__and3b_1
XFILLER_125_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10408_ _03535_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__clkbuf_1
X_14176_ _06911_ _06912_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__and2_1
XFILLER_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11388_ _04147_ gpout0.hpos\[2\] gpout0.hpos\[3\] _04162_ _04167_ vssd1 vssd1 vccd1
+ vccd1 _04168_ sky130_fd_sc_hd__o221a_1
XFILLER_125_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _03499_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_152_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13127_ _05859_ _05863_ _05811_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__mux2_1
XFILLER_140_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _02622_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__clkbuf_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17935_ _10110_ _09977_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__nor2_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _05759_ _05772_ _05775_ _05699_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__nor4b_2
XFILLER_100_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12009_ rbzero.tex_b1\[59\] rbzero.tex_b1\[58\] _04350_ vssd1 vssd1 vccd1 vccd1 _04784_
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17866_ _01561_ _01562_ _01568_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16817_ rbzero.debug_overlay.playerY\[-3\] vssd1 vssd1 vccd1 vccd1 _09459_ sky130_fd_sc_hd__clkinv_2
XFILLER_54_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17797_ _10239_ _08057_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__nor2_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19536_ _03010_ _03011_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__xnor2_1
X_16748_ _09245_ _08059_ _09389_ vssd1 vssd1 vccd1 vccd1 _09390_ sky130_fd_sc_hd__or3_1
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20165__192 clknet_1_0__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__inv_2
XFILLER_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19467_ _02904_ rbzero.wall_tracer.rayAddendY\[5\] vssd1 vssd1 vccd1 vccd1 _02948_
+ sky130_fd_sc_hd__nand2_1
XFILLER_146_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16679_ _09181_ _09158_ vssd1 vssd1 vccd1 vccd1 _09322_ sky130_fd_sc_hd__or2b_1
XFILLER_50_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18418_ _01928_ _02004_ _02003_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19398_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.debug_overlay.vplaneY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__and2_1
XFILLER_194_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18349_ _10248_ _09991_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__nor2_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21360_ net281 _01129_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21291_ clknet_leaf_37_i_clk _01060_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[9\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_6_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10690_ rbzero.tex_g1\[12\] rbzero.tex_g1\[13\] _03680_ vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21627_ clknet_leaf_28_i_clk _01396_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_201_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12360_ _05127_ _05099_ _05107_ net1 vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21558_ net479 _01327_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ _04075_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__or2_1
XFILLER_138_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20509_ _09750_ _03404_ _03405_ _03250_ rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1
+ _01399_ sky130_fd_sc_hd__a32o_1
X_12291_ _05042_ _05054_ _05059_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a21o_1
XFILLER_193_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21489_ net410 _01258_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14030_ _06762_ _06764_ _06765_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a21o_1
X_11242_ _04004_ _04022_ _04024_ _04025_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__and4b_2
XFILLER_84_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11173_ rbzero.othery\[2\] _03933_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__xnor2_1
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15981_ _07923_ vssd1 vssd1 vccd1 vccd1 _08626_ sky130_fd_sc_hd__inv_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17720_ _10195_ _10284_ vssd1 vssd1 vccd1 vccd1 _10285_ sky130_fd_sc_hd__xnor2_1
XFILLER_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14932_ rbzero.wall_tracer.visualWallDist\[2\] _07618_ vssd1 vssd1 vccd1 vccd1 _07631_
+ sky130_fd_sc_hd__or2_1
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20307__320 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__inv_2
X_17651_ _10095_ _10097_ _10093_ vssd1 vssd1 vccd1 vccd1 _10216_ sky130_fd_sc_hd__a21bo_1
X_14863_ rbzero.wall_tracer.stepDistY\[8\] _07579_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07580_ sky130_fd_sc_hd__mux2_1
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16602_ _07938_ vssd1 vssd1 vccd1 vccd1 _09245_ sky130_fd_sc_hd__buf_2
X_13814_ _06423_ _06550_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__xor2_1
X_17582_ _09994_ _10002_ vssd1 vssd1 vccd1 vccd1 _10148_ sky130_fd_sc_hd__nand2_1
XFILLER_17_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14794_ _00004_ _07524_ _07525_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__a21oi_1
XFILLER_91_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19321_ rbzero.spi_registers.new_vshift\[3\] rbzero.spi_registers.spi_buffer\[3\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__mux2_1
XFILLER_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16533_ _09175_ _09176_ vssd1 vssd1 vccd1 vccd1 _09177_ sky130_fd_sc_hd__xor2_1
XFILLER_17_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13745_ _06471_ _06472_ _06481_ _06474_ _06480_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__a32o_1
XFILLER_17_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10957_ rbzero.tex_b1\[13\] rbzero.tex_b1\[14\] _03817_ vssd1 vssd1 vccd1 vccd1 _03826_
+ sky130_fd_sc_hd__mux2_1
XFILLER_189_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19252_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_sky\[4\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__mux2_1
XFILLER_71_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16464_ _09106_ _09107_ vssd1 vssd1 vccd1 vccd1 _09108_ sky130_fd_sc_hd__nor2_1
XFILLER_204_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13676_ _06398_ _06412_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__xor2_1
XFILLER_143_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10888_ rbzero.tex_b1\[46\] rbzero.tex_b1\[47\] _03784_ vssd1 vssd1 vccd1 vccd1 _03790_
+ sky130_fd_sc_hd__mux2_1
X_18203_ _01802_ _01803_ _01901_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__and3_1
XFILLER_188_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15415_ rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendX\[-3\] rbzero.wall_tracer.side
+ vssd1 vssd1 vccd1 vccd1 _08060_ sky130_fd_sc_hd__mux2_1
XFILLER_176_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12627_ _05380_ vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__clkbuf_1
X_19183_ rbzero.floor_leak\[2\] _02732_ _02736_ _02722_ vssd1 vssd1 vccd1 vccd1 _00742_
+ sky130_fd_sc_hd__o211a_1
X_16395_ _09031_ _09039_ vssd1 vssd1 vccd1 vccd1 _09040_ sky130_fd_sc_hd__xnor2_2
X_18134_ _01833_ _01834_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__and2_1
XFILLER_185_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15346_ _05345_ _05466_ _07893_ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__mux2_1
XFILLER_200_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] _05300_
+ _05310_ _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a221o_1
XFILLER_106_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18065_ _01764_ _01765_ _01646_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11509_ _04210_ _04284_ _04288_ _04242_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__a211o_1
X_20353__362 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__inv_2
XFILLER_89_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15277_ _07916_ _07921_ vssd1 vssd1 vccd1 vccd1 _07922_ sky130_fd_sc_hd__or2_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12489_ rbzero.wall_tracer.trackDistY\[-11\] _05242_ rbzero.wall_tracer.trackDistY\[-12\]
+ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__o211a_1
XFILLER_144_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17016_ _09654_ _09655_ vssd1 vssd1 vccd1 vccd1 _09656_ sky130_fd_sc_hd__nand2_1
X_14228_ _06935_ _06963_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__or2_1
XFILLER_171_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ _06864_ _06895_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__xor2_1
XFILLER_4_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18967_ _02613_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__clkbuf_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17918_ _01498_ _01620_ _01618_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__o21ai_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18898_ rbzero.spi_registers.spi_counter\[0\] _02564_ _02567_ vssd1 vssd1 vccd1 vccd1
+ _02568_ sky130_fd_sc_hd__a21oi_1
XFILLER_152_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17849_ _05532_ _01552_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__nand2_1
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20860_ clknet_leaf_0_i_clk _00629_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19519_ _02983_ _02987_ _02996_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__nand3_1
X_20791_ clknet_leaf_29_i_clk _00560_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21412_ net333 _01181_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21343_ net264 _01112_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21274_ clknet_leaf_89_i_clk _01043_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20181__207 clknet_1_0__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__inv_2
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ rbzero.tex_g1\[5\] rbzero.tex_g1\[4\] _04336_ vssd1 vssd1 vccd1 vccd1 _04637_
+ sky130_fd_sc_hd__mux2_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10811_ _03749_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__clkbuf_1
X_11791_ rbzero.tex_g0\[55\] _04347_ _04348_ _04217_ vssd1 vssd1 vccd1 vccd1 _04569_
+ sky130_fd_sc_hd__a31o_1
XFILLER_14_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20989_ clknet_leaf_14_i_clk _00758_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13530_ _06219_ _06266_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__xor2_1
X_10742_ rbzero.tex_g0\[52\] rbzero.tex_g0\[51\] _03706_ vssd1 vssd1 vccd1 vccd1 _03713_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10673_ rbzero.tex_g1\[20\] rbzero.tex_g1\[21\] _03669_ vssd1 vssd1 vccd1 vccd1 _03677_
+ sky130_fd_sc_hd__mux2_1
X_13461_ _06172_ _06187_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__and2b_1
XFILLER_199_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15200_ _07851_ _07852_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__nand2_1
XFILLER_199_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12412_ _05146_ _04666_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__nand2_1
XFILLER_51_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16180_ _08822_ _08824_ vssd1 vssd1 vccd1 vccd1 _08825_ sky130_fd_sc_hd__nand2_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13392_ _06111_ _06128_ _06109_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__a21o_1
XFILLER_194_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15131_ _07783_ _07784_ _07786_ _07787_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__o211a_1
X_12343_ _04323_ _05084_ _05107_ net68 vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__a22oi_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12274_ _05032_ net20 vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__and2_1
X_15062_ _07710_ _07714_ _07711_ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__o21ai_1
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11225_ gpout0.hpos\[7\] vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__inv_2
X_14013_ _06748_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__nand2_1
XFILLER_49_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19870_ rbzero.debug_overlay.playerX\[3\] _03176_ vssd1 vssd1 vccd1 vccd1 _03180_
+ sky130_fd_sc_hd__nor2_1
XFILLER_150_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03039_ clknet_0__03039_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03039_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11156_ rbzero.debug_overlay.playerX\[4\] rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1
+ vccd1 _03945_ sky130_fd_sc_hd__xor2_1
X_18821_ _02499_ _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18752_ _02398_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__buf_6
X_15964_ _08586_ _08608_ vssd1 vssd1 vccd1 vccd1 _08609_ sky130_fd_sc_hd__xor2_1
XFILLER_23_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11087_ rbzero.tex_b0\[16\] rbzero.tex_b0\[15\] _03887_ vssd1 vssd1 vccd1 vccd1 _03894_
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17703_ _10130_ _10266_ _10267_ vssd1 vssd1 vccd1 vccd1 _10268_ sky130_fd_sc_hd__o21a_1
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14915_ rbzero.wall_tracer.visualWallDist\[-3\] _07618_ vssd1 vssd1 vccd1 vccd1 _07619_
+ sky130_fd_sc_hd__or2_1
X_18683_ _02235_ _02249_ _02378_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a21oi_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15895_ _08487_ _08506_ _08508_ vssd1 vssd1 vccd1 vccd1 _08540_ sky130_fd_sc_hd__and3_1
XFILLER_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ _10090_ _10108_ _10198_ vssd1 vssd1 vccd1 vccd1 _10199_ sky130_fd_sc_hd__a21o_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ rbzero.wall_tracer.stepDistY\[4\] _07566_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07567_ sky130_fd_sc_hd__mux2_1
XFILLER_63_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17565_ _08872_ _08873_ vssd1 vssd1 vccd1 vccd1 _10131_ sky130_fd_sc_hd__nand2_1
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14777_ _07473_ _07507_ _07509_ _05814_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__o211ai_1
XFILLER_95_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11989_ rbzero.tex_b1\[7\] rbzero.tex_b1\[6\] _04212_ vssd1 vssd1 vccd1 vccd1 _04764_
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19304_ rbzero.spi_registers.new_other\[7\] rbzero.spi_registers.spi_buffer\[7\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__mux2_1
XFILLER_189_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16516_ _09002_ _09019_ _09159_ vssd1 vssd1 vccd1 vccd1 _09160_ sky130_fd_sc_hd__a21bo_1
XFILLER_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13728_ _06436_ _06459_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__xor2_1
XFILLER_56_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17496_ _10060_ _10061_ vssd1 vssd1 vccd1 vccd1 _10062_ sky130_fd_sc_hd__xor2_1
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19235_ rbzero.spi_registers.new_vshift\[4\] _02763_ vssd1 vssd1 vccd1 vccd1 _02769_
+ sky130_fd_sc_hd__or2_1
X_16447_ _08961_ _08966_ vssd1 vssd1 vccd1 vccd1 _09091_ sky130_fd_sc_hd__nand2_1
X_13659_ _06381_ _06386_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_71_i_clk clknet_3_5_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_158_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19166_ rbzero.othery\[3\] _02710_ _02724_ _02722_ vssd1 vssd1 vccd1 vccd1 _00737_
+ sky130_fd_sc_hd__o211a_1
X_20277__293 clknet_1_0__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__inv_2
X_16378_ _08297_ _08326_ vssd1 vssd1 vccd1 vccd1 _09023_ sky130_fd_sc_hd__nor2_1
XFILLER_185_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18117_ _01728_ _01729_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__nor2_1
XFILLER_8_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15329_ _07970_ _07549_ _07973_ vssd1 vssd1 vccd1 vccd1 _07974_ sky130_fd_sc_hd__o21ai_4
X_19097_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.spi_buffer\[3\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__mux2_1
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18048_ _01748_ _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__xor2_1
XFILLER_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_86_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_67_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20010_ _04890_ _04989_ _02703_ _04990_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__or4b_1
XFILLER_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19999_ rbzero.pov.ready_buffer\[3\] _03246_ _03248_ rbzero.debug_overlay.vplaneY\[-6\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__a221o_1
XFILLER_154_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20912_ clknet_leaf_20_i_clk _00681_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ clknet_leaf_61_i_clk _00612_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20774_ clknet_leaf_39_i_clk _00543_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_1_0_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21326_ net247 _01095_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21257_ clknet_leaf_96_i_clk _01026_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_11_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11010_ _03853_ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21188_ clknet_leaf_26_i_clk _00957_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12961_ _05697_ _05692_ _05648_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__or3_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _05741_ _07397_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__nand2_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11912_ rbzero.tex_b0\[23\] rbzero.tex_b0\[22\] _04271_ vssd1 vssd1 vccd1 vccd1 _04688_
+ sky130_fd_sc_hd__mux2_1
X_15680_ _08298_ _08312_ vssd1 vssd1 vccd1 vccd1 _08325_ sky130_fd_sc_hd__nor2_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ rbzero.wall_tracer.visualWallDist\[3\] _04030_ vssd1 vssd1 vccd1 vccd1 _05629_
+ sky130_fd_sc_hd__nor2_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _07314_ _07367_ _07311_ _07313_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__o211ai_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _04379_ _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__or2_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _09915_ _09916_ vssd1 vssd1 vccd1 vccd1 _09917_ sky130_fd_sc_hd__nor2_2
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14562_ _07044_ _07089_ _07298_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__a21oi_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ rbzero.tex_g0\[30\] _04211_ _04125_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__a21o_1
XFILLER_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _08808_ _08810_ vssd1 vssd1 vccd1 vccd1 _08946_ sky130_fd_sc_hd__nor2_1
X_13513_ _06248_ _06249_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__nor2_1
X_10725_ rbzero.tex_g0\[60\] rbzero.tex_g0\[59\] _03624_ vssd1 vssd1 vccd1 vccd1 _03704_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17281_ rbzero.wall_tracer.trackDistX\[-6\] rbzero.wall_tracer.stepDistX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _09854_ sky130_fd_sc_hd__nor2_1
X_14493_ _07045_ _07046_ _07048_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__a21bo_1
X_19020_ _02641_ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16232_ _08194_ _08579_ vssd1 vssd1 vccd1 vccd1 _08877_ sky130_fd_sc_hd__or2_1
X_13444_ _05910_ _06176_ _06085_ _06180_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__a31oi_1
XFILLER_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10656_ rbzero.tex_g1\[28\] rbzero.tex_g1\[29\] _03658_ vssd1 vssd1 vccd1 vccd1 _03668_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16163_ _08666_ _08668_ vssd1 vssd1 vccd1 vccd1 _08808_ sky130_fd_sc_hd__xnor2_4
XFILLER_186_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10587_ _03631_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__clkbuf_1
X_13375_ _06061_ _05940_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__nor2_1
XFILLER_103_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15114_ _07758_ _07761_ _07771_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12326_ _05082_ net28 vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__and2_1
XFILLER_155_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16094_ _08695_ _08738_ vssd1 vssd1 vccd1 vccd1 _08739_ sky130_fd_sc_hd__xnor2_2
XFILLER_181_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15045_ rbzero.debug_overlay.vplaneX\[-7\] _07705_ vssd1 vssd1 vccd1 vccd1 _07708_
+ sky130_fd_sc_hd__or2_1
X_19922_ rbzero.debug_overlay.playerY\[0\] _03198_ _03219_ _03209_ vssd1 vssd1 vccd1
+ vccd1 _00998_ sky130_fd_sc_hd__o211a_1
X_12257_ _05021_ net64 _05024_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__a211o_1
XFILLER_69_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ _03987_ _03996_ _03955_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__o21a_1
X_12188_ _04666_ _04903_ _04904_ _04905_ _04958_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a41o_2
X_19853_ rbzero.debug_overlay.playerX\[-1\] _03139_ _03166_ net60 vssd1 vssd1 vccd1
+ vccd1 _00982_ sky130_fd_sc_hd__a211o_1
XFILLER_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18804_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.stepDistY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__or2_1
X_11139_ rbzero.debug_overlay.playerX\[1\] _03924_ _03925_ rbzero.debug_overlay.playerY\[0\]
+ _03927_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__a221o_1
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16996_ _09626_ _09635_ vssd1 vssd1 vccd1 vccd1 _09636_ sky130_fd_sc_hd__nand2_1
X_19784_ rbzero.pov.spi_buffer\[65\] rbzero.pov.spi_buffer\[66\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03121_ sky130_fd_sc_hd__mux2_1
XFILLER_84_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18735_ _09863_ _02424_ _02425_ _09843_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__o31ai_1
XFILLER_83_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15947_ _07601_ _04014_ _07990_ _07927_ vssd1 vssd1 vccd1 vccd1 _08592_ sky130_fd_sc_hd__and4_1
XFILLER_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18666_ _02353_ _02361_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__xnor2_1
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15878_ _08445_ _08250_ vssd1 vssd1 vccd1 vccd1 _08523_ sky130_fd_sc_hd__nand2_1
XFILLER_63_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14829_ _07527_ _07504_ _07449_ _07459_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_92_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17617_ _10179_ _10180_ _10175_ _10177_ vssd1 vssd1 vccd1 vccd1 _10182_ sky130_fd_sc_hd__o211a_1
X_18597_ _02169_ _02170_ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__or2b_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17548_ _09117_ _09693_ _09992_ _10113_ vssd1 vssd1 vccd1 vccd1 _10114_ sky130_fd_sc_hd__o31a_1
XFILLER_177_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17479_ _09952_ _10040_ _10044_ vssd1 vssd1 vccd1 vccd1 _10045_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19218_ rbzero.spi_registers.new_floor\[4\] rbzero.color_floor\[4\] _02751_ vssd1
+ vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__mux2_1
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20490_ rbzero.traced_texa\[1\] rbzero.texV\[1\] vssd1 vssd1 vccd1 vccd1 _03389_
+ sky130_fd_sc_hd__or2_1
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19149_ rbzero.spi_registers.new_other\[7\] _02712_ vssd1 vssd1 vccd1 vccd1 _02715_
+ sky130_fd_sc_hd__or2_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21111_ net201 _00880_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21042_ clknet_leaf_76_i_clk _00811_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ clknet_leaf_50_i_clk _00595_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_20293__308 clknet_1_1__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__inv_2
XFILLER_168_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20757_ clknet_leaf_36_i_clk _00526_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_126_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10510_ _03557_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__clkbuf_4
X_11490_ _04207_ _04233_ _04243_ _04269_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__a31o_1
XFILLER_156_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20688_ clknet_leaf_54_i_clk _00472_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10441_ rbzero.tex_r1\[0\] rbzero.tex_r1\[1\] _03549_ vssd1 vssd1 vccd1 vccd1 _03553_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10372_ rbzero.tex_r1\[33\] rbzero.tex_r1\[34\] _03516_ vssd1 vssd1 vccd1 vccd1 _03517_
+ sky130_fd_sc_hd__mux2_1
X_13160_ _05811_ _05819_ _05814_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a21o_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12111_ gpout0.vpos\[2\] vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__buf_2
XFILLER_108_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13091_ _05826_ _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__and2_1
X_21309_ net230 _01078_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12042_ _04813_ _04809_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__nor2_1
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16850_ _09489_ _09490_ vssd1 vssd1 vccd1 vccd1 _09491_ sky130_fd_sc_hd__and2b_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15801_ _08445_ _08227_ vssd1 vssd1 vccd1 vccd1 _08446_ sky130_fd_sc_hd__nand2_1
X_16781_ _09418_ _09422_ vssd1 vssd1 vccd1 vccd1 _09423_ sky130_fd_sc_hd__and2_1
X_13993_ _06724_ _06690_ _06728_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__o21bai_1
XFILLER_92_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18520_ _02215_ _02217_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__xnor2_2
XFILLER_207_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _08376_ vssd1 vssd1 vccd1 vccd1 _08377_ sky130_fd_sc_hd__buf_4
XFILLER_206_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ _05678_ _05679_ _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__mux2_1
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _02147_ _02148_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__xor2_2
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15663_ _08265_ _08307_ vssd1 vssd1 vccd1 vccd1 _08308_ sky130_fd_sc_hd__xnor2_1
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _04030_ _05338_ _05339_ _05611_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a31o_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _09967_ _09968_ vssd1 vssd1 vccd1 vccd1 _09969_ sky130_fd_sc_hd__xor2_2
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14614_ _05793_ _07350_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__and2_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _02070_ _02080_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__nand2_1
X_11826_ rbzero.tex_g1\[61\] rbzero.tex_g1\[60\] _04392_ vssd1 vssd1 vccd1 vccd1 _04603_
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15594_ _08238_ vssd1 vssd1 vccd1 vccd1 _08239_ sky130_fd_sc_hd__clkbuf_4
XFILLER_18_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _09898_ _09899_ _09900_ _09893_ vssd1 vssd1 vccd1 vccd1 _09901_ sky130_fd_sc_hd__o211ai_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _07276_ _07280_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__nor2_1
XFILLER_183_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11757_ rbzero.tex_g0\[2\] _04211_ _04125_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__a21o_1
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10708_ _03695_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__clkbuf_1
X_17264_ rbzero.wall_tracer.trackDistX\[-8\] rbzero.wall_tracer.stepDistX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _09839_ sky130_fd_sc_hd__and2_1
XFILLER_202_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14476_ _07211_ _07212_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__nor2_1
X_11688_ rbzero.debug_overlay.vplaneX\[-1\] _04465_ _04466_ rbzero.debug_overlay.vplaneX\[-8\]
+ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__a22o_1
X_19003_ _02632_ vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__clkbuf_1
X_16215_ _08858_ _08859_ vssd1 vssd1 vccd1 vccd1 _08860_ sky130_fd_sc_hd__xor2_1
X_13427_ _05991_ _05978_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__nor2_1
X_10639_ _03659_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__clkbuf_1
X_17195_ _05413_ vssd1 vssd1 vccd1 vccd1 _09780_ sky130_fd_sc_hd__inv_2
XFILLER_10_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16146_ _08782_ _08783_ _08786_ vssd1 vssd1 vccd1 vccd1 _08791_ sky130_fd_sc_hd__or3_1
XFILLER_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13358_ _05920_ _05975_ _06093_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__or3b_1
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12309_ _05034_ _05027_ _05069_ _05077_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__a31o_2
XFILLER_170_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16077_ _08008_ _08042_ vssd1 vssd1 vccd1 vccd1 _08722_ sky130_fd_sc_hd__nor2_1
X_13289_ _05946_ _05973_ _06007_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__or3_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15028_ _07683_ _07691_ _07692_ vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__a21boi_1
X_19905_ _07954_ _03141_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__nor2_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19836_ rbzero.pov.ready_buffer\[63\] _07914_ _03146_ vssd1 vssd1 vccd1 vccd1 _03154_
+ sky130_fd_sc_hd__mux2_1
XFILLER_96_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19767_ rbzero.pov.spi_buffer\[57\] rbzero.pov.spi_buffer\[58\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03112_ sky130_fd_sc_hd__mux2_1
X_16979_ _09537_ _09518_ vssd1 vssd1 vccd1 vccd1 _09619_ sky130_fd_sc_hd__or2b_1
Xinput3 i_gpout0_sel[1] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_8
XFILLER_37_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18718_ _02408_ _02409_ _02407_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__o21a_1
X_19698_ rbzero.pov.spi_buffer\[24\] rbzero.pov.spi_buffer\[25\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux2_1
XFILLER_149_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18649_ _02241_ _02245_ _02344_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_0__03298_ _03298_ vssd1 vssd1 vccd1 vccd1 clknet_0__03298_ sky130_fd_sc_hd__clkbuf_16
XFILLER_25_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21660_ clknet_leaf_79_i_clk _01429_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20611_ gpout4.clk_div\[1\] gpout4.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__nand2_1
X_21591_ net132 _01360_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20542_ _03430_ _03431_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__a21o_1
XFILLER_178_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20473_ _03367_ _03369_ _03368_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__a21boi_1
XFILLER_119_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20136__167 clknet_1_0__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__inv_2
XFILLER_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21025_ clknet_leaf_4_i_clk _00794_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10990_ _03717_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__clkbuf_4
XFILLER_56_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20301__315 clknet_1_1__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__inv_2
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _05409_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _04387_ _04388_ _04389_ _04226_ _04306_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__o221a_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ clknet_leaf_54_i_clk _00578_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12591_ _05337_ _05344_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__and2_1
XFILLER_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14330_ _07061_ _07066_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__xor2_1
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11542_ gpout0.vpos\[8\] gpout0.vpos\[7\] gpout0.vpos\[6\] vssd1 vssd1 vccd1 vccd1
+ _04322_ sky130_fd_sc_hd__and3_1
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ _06997_ _06725_ vssd1 vssd1 vccd1 vccd1 _06998_ sky130_fd_sc_hd__xnor2_1
X_11473_ _04123_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__clkbuf_8
X_16000_ _07994_ _08594_ vssd1 vssd1 vccd1 vccd1 _08645_ sky130_fd_sc_hd__nor2_1
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13212_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__clkbuf_2
X_10424_ rbzero.tex_r1\[8\] rbzero.tex_r1\[9\] _03538_ vssd1 vssd1 vccd1 vccd1 _03544_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14192_ _06805_ _06667_ _06928_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__or3b_1
XFILLER_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13143_ _05837_ _05841_ _05807_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__mux2_1
X_10355_ rbzero.tex_r1\[41\] rbzero.tex_r1\[42\] _03505_ vssd1 vssd1 vccd1 vccd1 _03508_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17951_ _01513_ _01533_ _01532_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__a21oi_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__buf_2
XFILLER_183_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16902_ _08242_ _09129_ _08283_ vssd1 vssd1 vccd1 vccd1 _09543_ sky130_fd_sc_hd__a21oi_1
X_12025_ rbzero.tex_b1\[39\] rbzero.tex_b1\[38\] _04250_ vssd1 vssd1 vccd1 vccd1 _04800_
+ sky130_fd_sc_hd__mux2_1
XFILLER_111_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17882_ _09526_ _09359_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__nor2_1
X_16833_ _09379_ _09471_ _09473_ vssd1 vssd1 vccd1 vccd1 _09474_ sky130_fd_sc_hd__a21oi_2
XFILLER_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16764_ _09114_ _08204_ _09271_ vssd1 vssd1 vccd1 vccd1 _09406_ sky130_fd_sc_hd__or3_1
X_19552_ rbzero.pov.spi_counter\[2\] rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\]
+ _03024_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__and4bb_1
XFILLER_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13976_ _05982_ _06663_ _06712_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__or3_1
XFILLER_207_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18503_ _02060_ _02101_ _02058_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a21oi_1
XFILLER_185_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15715_ _07931_ _08109_ vssd1 vssd1 vccd1 vccd1 _08360_ sky130_fd_sc_hd__nor2_1
X_12927_ _05660_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__inv_2
XFILLER_206_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16695_ _09336_ _09337_ vssd1 vssd1 vccd1 vccd1 _09338_ sky130_fd_sc_hd__xnor2_1
X_19483_ _02905_ _04471_ _02961_ _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__o22ai_1
XFILLER_206_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15646_ _07912_ _08276_ vssd1 vssd1 vccd1 vccd1 _08291_ sky130_fd_sc_hd__nor2_1
X_18434_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.stepDistX\[8\] vssd1
+ vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__and2_1
X_12858_ rbzero.wall_tracer.visualWallDist\[-9\] _05355_ rbzero.wall_tracer.rcp_sel\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__mux2_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18365_ _01996_ _01979_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__or2b_1
XFILLER_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11809_ _04585_ _04586_ _04217_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__mux2_1
XFILLER_15_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15577_ _07894_ _05494_ vssd1 vssd1 vccd1 vccd1 _08222_ sky130_fd_sc_hd__nand2_1
X_12789_ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__buf_6
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17316_ _09863_ _09883_ _09884_ _09885_ vssd1 vssd1 vccd1 vccd1 _09886_ sky130_fd_sc_hd__o31ai_1
XFILLER_193_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14528_ _07261_ _07263_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__nand2_1
X_18296_ _01981_ _01995_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__xor2_1
XFILLER_119_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17247_ _09821_ _09822_ _09823_ vssd1 vssd1 vccd1 vccd1 _09824_ sky130_fd_sc_hd__a21oi_1
XFILLER_179_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14459_ _07168_ _07183_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__or2b_1
XFILLER_127_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17178_ rbzero.traced_texa\[6\] _09770_ _09769_ rbzero.wall_tracer.visualWallDist\[6\]
+ vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__a22o_1
XFILLER_127_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16129_ _08772_ _08773_ vssd1 vssd1 vccd1 vccd1 _08774_ sky130_fd_sc_hd__or2b_1
XFILLER_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19819_ _02822_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03319_ clknet_0__03319_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03319_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21643_ clknet_leaf_31_i_clk _01412_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21574_ net495 _01343_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_41 net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_52 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20525_ _03411_ _03414_ _03412_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__a21boi_1
XANTENNA_74 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20456_ _03357_ _03358_ _03359_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a21o_1
XFILLER_197_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21008_ clknet_leaf_3_i_clk _00777_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20055__93 clknet_1_1__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__inv_2
X_13830_ _06565_ _06566_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__nand2_1
XFILLER_63_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13761_ _06462_ _06496_ _06426_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__a21bo_1
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10973_ _03834_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15500_ _08137_ _08143_ _08144_ vssd1 vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__a21o_1
X_12712_ _05439_ _05441_ _05418_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__a21bo_1
X_16480_ _09118_ _09123_ vssd1 vssd1 vccd1 vccd1 _09124_ sky130_fd_sc_hd__xnor2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _06384_ _06385_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15431_ _08074_ _08075_ _07965_ vssd1 vssd1 vccd1 vccd1 _08076_ sky130_fd_sc_hd__or3_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12643_ rbzero.debug_overlay.playerY\[3\] _05393_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05395_ sky130_fd_sc_hd__mux2_1
X_18150_ _01848_ _01849_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__and2_1
XFILLER_157_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15362_ rbzero.wall_tracer.visualWallDist\[-7\] _04014_ _05207_ vssd1 vssd1 vccd1
+ vccd1 _08007_ sky130_fd_sc_hd__a21oi_1
X_12574_ _05326_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__and2_1
X_17101_ _09082_ _09740_ vssd1 vssd1 vccd1 vccd1 _09741_ sky130_fd_sc_hd__xnor2_2
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14313_ _07048_ _07049_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18081_ _01572_ _01659_ _01782_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a21boi_1
XFILLER_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ rbzero.tex_r0\[30\] _04273_ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__a21o_1
X_15293_ _04013_ _07936_ _07937_ vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__a21oi_4
XFILLER_157_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17032_ _09545_ _09670_ _09671_ vssd1 vssd1 vccd1 vccd1 _09672_ sky130_fd_sc_hd__a21oi_2
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14244_ _06946_ _06961_ _06980_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__a21oi_1
X_11456_ _04234_ _04235_ _04226_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__mux2_1
XFILLER_125_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20119__151 clknet_1_0__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__inv_2
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ rbzero.tex_r1\[16\] rbzero.tex_r1\[17\] _03527_ vssd1 vssd1 vccd1 vccd1 _03535_
+ sky130_fd_sc_hd__mux2_1
XFILLER_109_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14175_ _06886_ _06910_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__nand2_1
X_11387_ _04147_ gpout0.hpos\[2\] _04163_ _04164_ _04166_ vssd1 vssd1 vccd1 vccd1
+ _04167_ sky130_fd_sc_hd__a221o_1
XFILLER_125_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13126_ _05861_ _05862_ _05807_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__mux2_1
X_10338_ rbzero.tex_r1\[49\] rbzero.tex_r1\[50\] _03494_ vssd1 vssd1 vccd1 vccd1 _03499_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ rbzero.pov.spi_buffer\[24\] rbzero.pov.ready_buffer\[24\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02622_ sky130_fd_sc_hd__mux2_1
XFILLER_112_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17934_ _08895_ _10139_ _08626_ _09989_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_26_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _05700_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__inv_2
XFILLER_94_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ rbzero.tex_b1\[56\] _04291_ _04139_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a21o_1
XFILLER_61_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17865_ _01566_ _01567_ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__nand2_1
XFILLER_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xnet99_2 clknet_1_1__leaf__04835_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__inv_2
XFILLER_94_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19604_ clknet_1_0__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__buf_1
X_16816_ _09341_ _09457_ vssd1 vssd1 vccd1 vccd1 _09458_ sky130_fd_sc_hd__xnor2_4
XFILLER_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17796_ _01497_ _01499_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__nand2_1
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19535_ _02906_ rbzero.wall_tracer.rayAddendY\[10\] vssd1 vssd1 vccd1 vccd1 _03011_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16747_ _09387_ _09388_ vssd1 vssd1 vccd1 vccd1 _09389_ sky130_fd_sc_hd__nand2_1
X_13959_ _06080_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16678_ _09318_ _09320_ vssd1 vssd1 vccd1 vccd1 _09321_ sky130_fd_sc_hd__xnor2_1
X_19466_ rbzero.wall_tracer.rayAddendY\[4\] _00013_ _02947_ vssd1 vssd1 vccd1 vccd1
+ _00814_ sky130_fd_sc_hd__o21a_1
XFILLER_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18417_ _02105_ _02115_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__xnor2_2
X_15629_ _05193_ _08273_ _04013_ vssd1 vssd1 vccd1 vccd1 _08274_ sky130_fd_sc_hd__o21a_1
XFILLER_107_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19397_ _02865_ _02875_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__nand2_1
XFILLER_148_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18348_ _10266_ _02045_ _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__o21ba_1
XFILLER_148_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18279_ _01865_ _01873_ _01978_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a21o_1
XFILLER_174_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21290_ clknet_leaf_37_i_clk _01059_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[8\] sky130_fd_sc_hd__dfxtp_1
Xinput50 i_vec_csb vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_8
XFILLER_190_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20330__341 clknet_1_0__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__inv_2
XFILLER_131_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20172_ clknet_1_1__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__buf_1
XFILLER_104_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20248__268 clknet_1_0__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__inv_2
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19588__44 clknet_1_0__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__inv_2
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21626_ clknet_leaf_28_i_clk _01395_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21557_ net478 _01326_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _04071_ _04074_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__and2_1
X_20508_ _03401_ _03402_ _03403_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__nand3_1
X_12290_ _05055_ _05056_ _05057_ _05058_ _05033_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__o311a_1
XFILLER_193_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21488_ net409 _01257_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11241_ _03475_ _04006_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__nor2_1
XFILLER_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20439_ _03343_ _03344_ _03345_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__or3_1
XFILLER_101_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ rbzero.otherx\[4\] rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1 vccd1 _03961_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_84_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15980_ _07912_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08625_ sky130_fd_sc_hd__or3_1
XFILLER_121_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14931_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.trackDistX\[2\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__mux2_1
XFILLER_76_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17650_ _10073_ _10077_ _10075_ vssd1 vssd1 vccd1 vccd1 _10215_ sky130_fd_sc_hd__a21bo_1
XFILLER_76_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14862_ _07456_ _07577_ _07578_ _07487_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__o31a_2
XFILLER_75_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16601_ _07932_ _07938_ _08035_ _08046_ vssd1 vssd1 vccd1 vccd1 _09244_ sky130_fd_sc_hd__or4_1
X_13813_ _06426_ _06462_ _06422_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__o21bai_1
X_17581_ _10122_ _10146_ vssd1 vssd1 vccd1 vccd1 _10147_ sky130_fd_sc_hd__xnor2_2
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14793_ rbzero.wall_tracer.stepDistY\[-7\] _00004_ vssd1 vssd1 vccd1 vccd1 _07525_
+ sky130_fd_sc_hd__nor2_1
XFILLER_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16532_ _09031_ _09039_ _09037_ vssd1 vssd1 vccd1 vccd1 _09176_ sky130_fd_sc_hd__a21oi_2
X_19320_ _02816_ vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__clkbuf_1
X_13744_ _06474_ _06480_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__xor2_1
XFILLER_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10956_ _03825_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16463_ _09102_ _09105_ vssd1 vssd1 vccd1 vccd1 _09107_ sky130_fd_sc_hd__and2_1
X_19251_ _02778_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__clkbuf_1
X_13675_ _06405_ _06410_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__o21ba_1
X_10887_ _03789_ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__clkbuf_1
X_18202_ _01902_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__inv_2
X_15414_ _08058_ vssd1 vssd1 vccd1 vccd1 _08059_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12626_ _05379_ _03942_ _05284_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__mux2_1
X_19182_ rbzero.spi_registers.new_leak\[2\] _02733_ vssd1 vssd1 vccd1 vccd1 _02736_
+ sky130_fd_sc_hd__or2_1
X_16394_ _09037_ _09038_ vssd1 vssd1 vccd1 vccd1 _09039_ sky130_fd_sc_hd__nor2_1
X_18133_ _01831_ _01832_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__nand2_1
XFILLER_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15345_ _05196_ vssd1 vssd1 vccd1 vccd1 _07990_ sky130_fd_sc_hd__buf_4
X_12557_ rbzero.debug_overlay.facingY\[-2\] rbzero.wall_tracer.rayAddendY\[6\] rbzero.wall_tracer.rayAddendY\[5\]
+ rbzero.debug_overlay.facingY\[-3\] vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__o211a_1
XFILLER_89_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18064_ _01646_ _01764_ _01765_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__and3_1
X_11508_ _04285_ _04286_ _04287_ _04226_ _04230_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__o221a_1
X_15276_ _07920_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__clkinv_2
X_12488_ rbzero.wall_tracer.trackDistX\[-12\] vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__inv_2
XFILLER_176_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17015_ _09618_ _09619_ _09653_ vssd1 vssd1 vccd1 vccd1 _09655_ sky130_fd_sc_hd__nand3_1
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14227_ _06935_ _06963_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__nand2_1
XFILLER_172_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11439_ _04218_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__buf_4
XFILLER_144_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14158_ _06776_ _06677_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__nor2_1
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _05835_ _05845_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__nor2_4
XFILLER_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14089_ _06806_ _06808_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__xnor2_1
X_18966_ rbzero.pov.spi_buffer\[16\] rbzero.pov.ready_buffer\[16\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02613_ sky130_fd_sc_hd__mux2_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17917_ _08057_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__buf_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18897_ rbzero.spi_registers.spi_counter\[6\] rbzero.spi_registers.spi_counter\[5\]
+ rbzero.spi_registers.spi_counter\[4\] vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__or3_1
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17848_ _01550_ _01551_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__xnor2_2
XFILLER_94_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17779_ _01473_ _01481_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__or2_1
XFILLER_148_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19518_ rbzero.debug_overlay.vplaneY\[0\] _02980_ _02993_ _02995_ vssd1 vssd1 vccd1
+ vccd1 _02996_ sky130_fd_sc_hd__o22a_1
XFILLER_207_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20790_ clknet_leaf_47_i_clk _00559_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19449_ _02930_ _02931_ _02911_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__o21bai_1
XFILLER_195_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21411_ net332 _01180_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21342_ net263 _01111_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21273_ clknet_leaf_93_i_clk _01042_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_162_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ rbzero.tex_g0\[20\] rbzero.tex_g0\[19\] _03740_ vssd1 vssd1 vccd1 vccd1 _03749_
+ sky130_fd_sc_hd__mux2_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ rbzero.tex_g0\[54\] _04350_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__and2_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20988_ clknet_leaf_10_i_clk _00757_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_207_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10741_ _03712_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13460_ _06170_ _06171_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and2b_1
X_10672_ _03676_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12411_ _05150_ _05138_ _05152_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a31o_2
XFILLER_90_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21609_ net126 _01378_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13391_ _06126_ _06127_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__nor2_1
XFILLER_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15130_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[3\] vssd1
+ vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__or2_1
X_12342_ _05101_ _05105_ _05109_ net28 vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__o22a_1
XFILLER_194_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15061_ _07721_ _07722_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__nand2_1
X_12273_ net23 _05033_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__nor2_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14012_ _06746_ _06747_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__or2_1
X_11224_ _04010_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_4
XFILLER_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03038_ clknet_0__03038_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03038_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18820_ _02492_ _02494_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__or2_1
X_11155_ rbzero.debug_overlay.playerY\[1\] _03942_ vssd1 vssd1 vccd1 vccd1 _03944_
+ sky130_fd_sc_hd__or2_1
X_18751_ _09863_ _02438_ _02439_ _09860_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__o31ai_1
X_11086_ _03893_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15963_ _08605_ _08606_ _08607_ vssd1 vssd1 vccd1 vccd1 _08608_ sky130_fd_sc_hd__a21oi_1
XFILLER_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17702_ _10139_ _08873_ _08263_ _10134_ vssd1 vssd1 vccd1 vccd1 _10267_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14914_ _07594_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__clkbuf_2
X_18682_ _02250_ _02287_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__and2b_1
X_15894_ _08512_ _08538_ vssd1 vssd1 vccd1 vccd1 _08539_ sky130_fd_sc_hd__xor2_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ _10092_ _10107_ vssd1 vssd1 vccd1 vccd1 _10198_ sky130_fd_sc_hd__nor2_1
XFILLER_64_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14845_ _05929_ _07456_ _07458_ _07487_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__o31a_2
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17564_ _08872_ _08873_ _10129_ vssd1 vssd1 vccd1 vccd1 _10130_ sky130_fd_sc_hd__or3_1
X_14776_ _07477_ _07475_ _07508_ _05884_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__a211o_1
X_11988_ rbzero.tex_b1\[5\] rbzero.tex_b1\[4\] _04212_ vssd1 vssd1 vccd1 vccd1 _04763_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19303_ _02807_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16515_ _09020_ _09000_ vssd1 vssd1 vccd1 vccd1 _09159_ sky130_fd_sc_hd__or2b_1
X_13727_ _06423_ _06463_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__nand2_1
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10939_ _03816_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17495_ _09096_ _09217_ vssd1 vssd1 vccd1 vccd1 _10061_ sky130_fd_sc_hd__nor2_1
XFILLER_182_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19234_ rbzero.spi_registers.vshift\[3\] _02762_ _02768_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00761_ sky130_fd_sc_hd__o211a_1
X_16446_ _09008_ _09018_ _09016_ vssd1 vssd1 vccd1 vccd1 _09090_ sky130_fd_sc_hd__a21o_1
X_13658_ _06352_ _06367_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _05318_ _05308_ _05312_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__or3_1
X_16377_ _08998_ _09021_ vssd1 vssd1 vccd1 vccd1 _09022_ sky130_fd_sc_hd__xnor2_4
X_19165_ rbzero.spi_registers.new_other\[3\] _02712_ vssd1 vssd1 vccd1 vccd1 _02724_
+ sky130_fd_sc_hd__or2_1
XFILLER_158_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13589_ _06325_ _06301_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18116_ _01691_ _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__xnor2_1
XFILLER_8_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15328_ _07971_ _05340_ _07972_ _05193_ vssd1 vssd1 vccd1 vccd1 _07973_ sky130_fd_sc_hd__a211o_1
XFILLER_173_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19096_ _02681_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18047_ _01503_ _01623_ _01624_ _01625_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_172_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15259_ _07903_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__clkbuf_4
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19998_ rbzero.pov.ready_buffer\[2\] _03239_ _03242_ rbzero.debug_overlay.vplaneY\[-7\]
+ _03254_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__o221a_1
XFILLER_98_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18949_ rbzero.pov.spi_buffer\[8\] rbzero.pov.ready_buffer\[8\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02604_ sky130_fd_sc_hd__mux2_1
XFILLER_67_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20911_ clknet_leaf_78_i_clk _00680_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_67_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20842_ clknet_leaf_61_i_clk _00611_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20773_ clknet_leaf_39_i_clk _00542_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21325_ net246 _01094_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21256_ clknet_leaf_84_i_clk _01025_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_132_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21187_ clknet_leaf_74_i_clk _00956_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20138_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__buf_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12960_ _05615_ _05639_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__xnor2_2
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _04271_ vssd1 vssd1 vccd1 vccd1 _04687_
+ sky130_fd_sc_hd__mux2_1
XFILLER_100_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12891_ _05627_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__buf_2
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _07306_ _07307_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__and2_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ rbzero.tex_g1\[33\] rbzero.tex_g1\[32\] _04337_ vssd1 vssd1 vccd1 vccd1 _04619_
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _07086_ _07088_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__nor2_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ rbzero.tex_g0\[31\] _04135_ _04136_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__and3_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13512_ _06237_ _06238_ _06247_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__and3_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _08620_ _08670_ vssd1 vssd1 vccd1 vccd1 _08945_ sky130_fd_sc_hd__xnor2_1
XFILLER_202_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10724_ _03703_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17280_ _09853_ vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__clkbuf_1
X_14492_ _07165_ _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__xnor2_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ _08867_ _08875_ vssd1 vssd1 vccd1 vccd1 _08876_ sky130_fd_sc_hd__nand2_1
X_13443_ _06041_ _06080_ _06084_ _05990_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__o22a_1
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10655_ _03667_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16162_ _08801_ _08805_ _08806_ vssd1 vssd1 vccd1 vccd1 _08807_ sky130_fd_sc_hd__a21oi_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13374_ _06109_ _06110_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__nor2_1
XFILLER_177_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10586_ rbzero.tex_g1\[61\] rbzero.tex_g1\[62\] _03549_ vssd1 vssd1 vccd1 vccd1 _03631_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15113_ _07769_ _07770_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__nand2_1
XFILLER_86_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12325_ _05087_ net64 _05091_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a211o_1
XFILLER_103_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16093_ _08716_ _08715_ vssd1 vssd1 vccd1 vccd1 _08738_ sky130_fd_sc_hd__and2b_1
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15044_ rbzero.wall_tracer.rayAddendX\[-4\] _00013_ _07702_ _07707_ vssd1 vssd1 vccd1
+ vccd1 _00492_ sky130_fd_sc_hd__o22a_1
X_19921_ rbzero.pov.ready_buffer\[53\] _03141_ _03192_ _03218_ vssd1 vssd1 vccd1 vccd1
+ _03219_ sky130_fd_sc_hd__a211o_1
X_12256_ _05021_ _04738_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__nor2_1
XFILLER_177_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11207_ _03993_ _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__nand2_2
X_19852_ _08093_ _03164_ _03143_ _03165_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__a211oi_1
X_12187_ _04907_ _04908_ net13 _04917_ _04957_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__o41a_2
XFILLER_123_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18803_ _02485_ _10028_ rbzero.wall_tracer.trackDistY\[0\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00613_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_150_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11138_ rbzero.debug_overlay.playerY\[3\] _03921_ _03926_ rbzero.map_rom.f3 vssd1
+ vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__a2bb2o_1
X_19783_ _03120_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__clkbuf_1
X_16995_ _09633_ _09634_ vssd1 vssd1 vccd1 vccd1 _09635_ sky130_fd_sc_hd__and2_1
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18734_ _02421_ _02422_ _02423_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__o21a_1
XFILLER_49_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11069_ _03884_ vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__clkbuf_1
X_15946_ rbzero.wall_tracer.visualWallDist\[-11\] _04014_ _05197_ _07992_ vssd1 vssd1
+ vccd1 vccd1 _08591_ sky130_fd_sc_hd__and4_1
XFILLER_77_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18665_ _02359_ _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__xnor2_1
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15877_ _08520_ _08521_ vssd1 vssd1 vccd1 vccd1 _08522_ sky130_fd_sc_hd__xnor2_1
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17616_ _10175_ _10177_ _10179_ _10180_ vssd1 vssd1 vccd1 vccd1 _10181_ sky130_fd_sc_hd__a211oi_1
XFILLER_63_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14828_ _00004_ _07552_ _07553_ vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__a21oi_1
X_18596_ _02166_ _02197_ _02292_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a21bo_1
XFILLER_64_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17547_ _08873_ _09991_ _09696_ vssd1 vssd1 vccd1 vccd1 _10113_ sky130_fd_sc_hd__or3b_1
X_14759_ _07357_ _07370_ vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__and2b_1
XFILLER_177_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17478_ _10042_ _10043_ vssd1 vssd1 vccd1 vccd1 _10044_ sky130_fd_sc_hd__or2_1
XFILLER_32_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19217_ rbzero.color_floor\[3\] _02751_ _02757_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__a21o_1
X_16429_ _09068_ _09072_ _09073_ vssd1 vssd1 vccd1 vccd1 _09074_ sky130_fd_sc_hd__a21o_1
XFILLER_146_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19148_ rbzero.otherx\[0\] _02710_ _02713_ _02714_ vssd1 vssd1 vccd1 vccd1 _00729_
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19079_ rbzero.pov.spi_buffer\[70\] rbzero.pov.ready_buffer\[70\] _02594_ vssd1 vssd1
+ vccd1 vccd1 _02672_ sky130_fd_sc_hd__mux2_1
XFILLER_106_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21110_ net200 _00879_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21041_ clknet_leaf_77_i_clk _00810_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20389__15 clknet_1_1__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__inv_2
XFILLER_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20825_ clknet_leaf_45_i_clk _00594_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20756_ clknet_leaf_40_i_clk _00525_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20687_ clknet_leaf_54_i_clk _00471_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10440_ _03552_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10371_ _03482_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__clkbuf_4
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ _04869_ _04879_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__nor2_1
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21308_ net229 _01077_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[15\] sky130_fd_sc_hd__dfxtp_1
X_13090_ _05591_ _05803_ _05796_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__mux2_1
XFILLER_152_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12041_ _04317_ _04814_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__or2_1
XFILLER_151_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21239_ clknet_leaf_68_i_clk _01008_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
X_20113__146 clknet_1_1__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__inv_2
Xclkbuf_opt_6_1_i_clk clknet_opt_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_6_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15800_ _07904_ rbzero.wall_tracer.stepDistY\[-1\] _08272_ _08274_ vssd1 vssd1 vccd1
+ vccd1 _08445_ sky130_fd_sc_hd__a22o_4
X_16780_ _09419_ _09421_ vssd1 vssd1 vccd1 vccd1 _09422_ sky130_fd_sc_hd__xnor2_1
X_13992_ _06724_ _06610_ _06728_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__or3b_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12943_ _05601_ _05638_ _05649_ _05628_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__o31a_1
X_15731_ _05206_ _08215_ vssd1 vssd1 vccd1 vccd1 _08376_ sky130_fd_sc_hd__or2_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _08356_ _09138_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__nor2_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15662_ _08276_ _07989_ vssd1 vssd1 vccd1 vccd1 _08307_ sky130_fd_sc_hd__nor2_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12874_ rbzero.wall_tracer.visualWallDist\[-2\] _05571_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05611_ sky130_fd_sc_hd__a21o_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _09545_ _09670_ _09672_ _09669_ vssd1 vssd1 vccd1 vccd1 _09968_ sky130_fd_sc_hd__a22oi_4
Xclkbuf_leaf_85_i_clk clknet_opt_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ rbzero.tex_g1\[63\] rbzero.tex_g1\[62\] _04337_ vssd1 vssd1 vccd1 vccd1 _04602_
+ sky130_fd_sc_hd__mux2_1
X_14613_ _07284_ _07321_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__xor2_1
XFILLER_92_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18381_ _02078_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__and2_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15593_ rbzero.wall_tracer.visualWallDist\[-12\] _04014_ vssd1 vssd1 vccd1 vccd1
+ _08238_ sky130_fd_sc_hd__nand2_4
XFILLER_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _07276_ _07280_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__and2_1
X_17332_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09900_ sky130_fd_sc_hd__nand2_1
XFILLER_57_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11756_ rbzero.tex_g0\[3\] _04088_ _04127_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__and3_1
XFILLER_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10707_ rbzero.tex_g1\[4\] rbzero.tex_g1\[5\] _03691_ vssd1 vssd1 vccd1 vccd1 _03695_
+ sky130_fd_sc_hd__mux2_1
XFILLER_186_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14475_ _07144_ _07156_ _07158_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__o21ba_1
X_17263_ rbzero.wall_tracer.trackDistX\[-8\] rbzero.wall_tracer.stepDistX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _09838_ sky130_fd_sc_hd__nor2_1
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11687_ _04437_ _04447_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__and2_2
X_19002_ rbzero.pov.spi_buffer\[33\] rbzero.pov.ready_buffer\[33\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02632_ sky130_fd_sc_hd__mux2_1
XFILLER_186_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16214_ _08816_ _08823_ vssd1 vssd1 vccd1 vccd1 _08859_ sky130_fd_sc_hd__nor2_1
X_13426_ _06160_ _06162_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__xor2_1
X_10638_ rbzero.tex_g1\[37\] rbzero.tex_g1\[38\] _03658_ vssd1 vssd1 vccd1 vccd1 _03659_
+ sky130_fd_sc_hd__mux2_1
X_17194_ _04019_ _05412_ vssd1 vssd1 vccd1 vccd1 _09779_ sky130_fd_sc_hd__nor2_4
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16145_ _08768_ _08789_ vssd1 vssd1 vccd1 vccd1 _08790_ sky130_fd_sc_hd__xnor2_1
X_13357_ _05991_ _05975_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__o21bai_1
X_10569_ rbzero.tex_r0\[6\] rbzero.tex_r0\[5\] _03613_ vssd1 vssd1 vccd1 vccd1 _03622_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12308_ _05072_ _05074_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__and3_1
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16076_ _08675_ _08720_ vssd1 vssd1 vccd1 vccd1 _08721_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_23_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13288_ _05983_ _06016_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__nor2_1
XFILLER_29_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15027_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__nand2_1
X_19904_ rbzero.debug_overlay.playerY\[-5\] _03198_ _03206_ _03157_ vssd1 vssd1 vccd1
+ vccd1 _00993_ sky130_fd_sc_hd__o211a_1
X_12239_ _05004_ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__nand2_1
XFILLER_170_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19835_ _03139_ _03152_ _03153_ _02765_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__o211a_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20088__123 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__inv_2
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_i_clk clknet_opt_9_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19766_ _03111_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16978_ _09536_ _09520_ vssd1 vssd1 vccd1 vccd1 _09618_ sky130_fd_sc_hd__or2b_1
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput4 i_gpout0_sel[2] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_8
XFILLER_83_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18717_ _02407_ _02408_ _02409_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__nor3_1
X_15929_ _08124_ _08490_ _08084_ vssd1 vssd1 vccd1 vccd1 _08574_ sky130_fd_sc_hd__a21oi_1
X_19697_ _03075_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18648_ _02045_ _02150_ _02152_ _02243_ _02343_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__a311o_1
Xclkbuf_0__03297_ _03297_ vssd1 vssd1 vccd1 vccd1 clknet_0__03297_ sky130_fd_sc_hd__clkbuf_16
XFILLER_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18579_ _01860_ _08423_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__nor2_1
XFILLER_149_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20610_ gpout4.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__nor2_1
XFILLER_33_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21590_ net131 _01359_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20541_ _03424_ _03428_ _03425_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__o21ai_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20472_ _03372_ _03373_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__or2_1
XFILLER_146_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21024_ clknet_leaf_94_i_clk _00793_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11610_ rbzero.tex_r1\[53\] rbzero.tex_r1\[52\] _04338_ vssd1 vssd1 vccd1 vccd1 _04389_
+ sky130_fd_sc_hd__mux2_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20808_ clknet_leaf_53_i_clk _00577_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12590_ _05309_ _05343_ _05305_ _05299_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__a211o_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11541_ gpout0.vpos\[3\] _04315_ _04316_ gpout0.vpos\[4\] _04320_ vssd1 vssd1 vccd1
+ vccd1 _04321_ sky130_fd_sc_hd__o221ai_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20739_ clknet_leaf_46_i_clk _00508_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.wall\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ _06134_ _06667_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__or2_1
XFILLER_183_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _04225_ _04251_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__or2_1
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ _05946_ _05947_ _05888_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__or3_1
XFILLER_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10423_ _03543_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14191_ _06895_ _06925_ _06927_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__a21oi_1
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13142_ _05830_ _05878_ _05778_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__mux2_2
X_10354_ _03507_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_174_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17950_ _01632_ _01652_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__xnor2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13073_ _05797_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__and2_1
XFILLER_151_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16901_ _09541_ vssd1 vssd1 vccd1 vccd1 _09542_ sky130_fd_sc_hd__inv_2
X_12024_ _04266_ _04798_ _04229_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__o21a_1
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17881_ _01581_ _01583_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__nand2_1
X_16832_ _09358_ _09360_ _09472_ vssd1 vssd1 vccd1 vccd1 _09473_ sky130_fd_sc_hd__o21a_1
XFILLER_116_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19551_ rbzero.pov.spi_counter\[5\] rbzero.pov.spi_counter\[4\] rbzero.pov.spi_counter\[3\]
+ rbzero.pov.spi_counter\[6\] vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__and4bb_1
XFILLER_47_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16763_ _09383_ _09404_ vssd1 vssd1 vccd1 vccd1 _09405_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13975_ _06659_ _06711_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18502_ _02163_ _02199_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15714_ _07940_ _08084_ vssd1 vssd1 vccd1 vccd1 _08359_ sky130_fd_sc_hd__nor2_1
XFILLER_47_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19482_ _02905_ rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1 _02962_
+ sky130_fd_sc_hd__and2_1
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ _05574_ _05662_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__xnor2_1
X_16694_ _09198_ _09200_ _09197_ vssd1 vssd1 vccd1 vccd1 _09337_ sky130_fd_sc_hd__a21o_1
XFILLER_73_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18433_ rbzero.wall_tracer.trackDistX\[8\] rbzero.wall_tracer.stepDistX\[8\] vssd1
+ vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__nor2_1
XFILLER_61_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15645_ _07977_ _07923_ vssd1 vssd1 vccd1 vccd1 _08290_ sky130_fd_sc_hd__nor2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _05589_ _05591_ _05593_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__or3_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18364_ _01995_ _01981_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__or2b_1
XFILLER_159_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11808_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _04341_ vssd1 vssd1 vccd1 vccd1 _04586_
+ sky130_fd_sc_hd__mux2_1
XFILLER_203_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15576_ _07566_ _08220_ _07970_ vssd1 vssd1 vccd1 vccd1 _08221_ sky130_fd_sc_hd__a21oi_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _04016_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__buf_4
XFILLER_187_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17315_ _09807_ _09458_ vssd1 vssd1 vccd1 vccd1 _09885_ sky130_fd_sc_hd__or2_1
XFILLER_109_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14527_ _07261_ _07263_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__nor2_1
X_11739_ _04320_ _04508_ _04517_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__and3_1
X_18295_ _01987_ _01994_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__xnor2_1
X_17246_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ _09815_ vssd1 vssd1 vccd1 vccd1 _09823_ sky130_fd_sc_hd__a21o_1
XFILLER_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14458_ _07162_ _07194_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__xnor2_1
XFILLER_179_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13409_ _06139_ _06140_ vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__nand2_1
X_14389_ _06698_ _07121_ _06760_ _07125_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__o31a_1
X_17177_ rbzero.traced_texa\[5\] _09770_ _09769_ rbzero.wall_tracer.visualWallDist\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a22o_1
XFILLER_143_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16128_ _08728_ _08731_ vssd1 vssd1 vccd1 vccd1 _08773_ sky130_fd_sc_hd__xnor2_1
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16059_ _08702_ _08703_ vssd1 vssd1 vccd1 vccd1 _08704_ sky130_fd_sc_hd__xor2_2
XFILLER_170_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19818_ rbzero.debug_overlay.playerX\[-9\] vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__inv_2
XFILLER_97_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03318_ clknet_0__03318_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03318_
+ sky130_fd_sc_hd__clkbuf_16
X_19749_ _03102_ vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21642_ clknet_leaf_32_i_clk _01411_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20142__172 clknet_1_1__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__inv_2
XFILLER_178_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_20 _09611_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21573_ net494 _01342_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_31 net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_42 _02406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20524_ _03416_ _03417_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__and2b_1
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_64 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_75 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20455_ _03357_ _03358_ _03359_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__nand3_1
XFILLER_180_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21007_ clknet_leaf_11_i_clk _00776_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13760_ _06426_ _06462_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__nand3b_1
XFILLER_44_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10972_ rbzero.tex_b1\[6\] rbzero.tex_b1\[7\] _03828_ vssd1 vssd1 vccd1 vccd1 _03834_
+ sky130_fd_sc_hd__mux2_1
X_20225__247 clknet_1_0__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__inv_2
XFILLER_189_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12711_ _05457_ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__xnor2_2
X_13691_ _05824_ _06134_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__or2_1
XFILLER_44_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15430_ _07964_ vssd1 vssd1 vccd1 vccd1 _08075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12642_ _05203_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__buf_4
XFILLER_54_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ _08002_ _08005_ vssd1 vssd1 vccd1 vccd1 _08006_ sky130_fd_sc_hd__nand2_1
XFILLER_106_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12573_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[11\] vssd1
+ vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__or2_1
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17100_ rbzero.debug_overlay.playerY\[-1\] rbzero.debug_overlay.playerX\[-1\] _07895_
+ vssd1 vssd1 vccd1 vccd1 _09740_ sky130_fd_sc_hd__mux2_1
X_11524_ _04217_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__buf_6
XFILLER_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14312_ _06724_ _06678_ _07047_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__o21bai_1
X_18080_ _01658_ _01656_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__or2b_1
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15292_ _07903_ rbzero.wall_tracer.stepDistY\[-5\] _05195_ vssd1 vssd1 vccd1 vccd1
+ _07937_ sky130_fd_sc_hd__a21o_1
XFILLER_178_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17031_ _07959_ _09276_ _08111_ _09126_ vssd1 vssd1 vccd1 vccd1 _09671_ sky130_fd_sc_hd__o22a_1
X_14243_ _06947_ _06948_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__xor2_1
X_11455_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _04214_ vssd1 vssd1 vccd1 vccd1 _04235_
+ sky130_fd_sc_hd__mux2_1
XFILLER_172_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10406_ _03534_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14174_ _06886_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__or2_1
XFILLER_178_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11386_ _04164_ gpout0.hpos\[1\] gpout0.hpos\[0\] _04165_ vssd1 vssd1 vccd1 vccd1
+ _04166_ sky130_fd_sc_hd__o211a_1
XFILLER_152_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13125_ _05728_ _05744_ _05791_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__mux2_1
X_10337_ _03498_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18982_ _02621_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _08767_ _10139_ _01518_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__or3b_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__clkbuf_4
XFILLER_97_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12007_ rbzero.tex_b1\[57\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__and3_1
X_17864_ _01563_ _01565_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__or2_1
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16815_ _09342_ _09456_ vssd1 vssd1 vccd1 vccd1 _09457_ sky130_fd_sc_hd__xor2_4
Xnet99_3 clknet_1_1__leaf__04835_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__inv_2
XFILLER_4_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17795_ _09276_ _08493_ _08044_ _01498_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__o22ai_1
XFILLER_66_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19534_ _02906_ rbzero.wall_tracer.rayAddendY\[9\] _03003_ vssd1 vssd1 vccd1 vccd1
+ _03010_ sky130_fd_sc_hd__a21oi_1
X_16746_ _07996_ _08129_ _08047_ _08705_ vssd1 vssd1 vccd1 vccd1 _09388_ sky130_fd_sc_hd__o22ai_1
XFILLER_81_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13958_ _06687_ _06694_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__or2_1
XFILLER_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19465_ _04035_ _02936_ _02937_ _02946_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a31o_1
X_12909_ _05610_ _05612_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__nand2_2
XFILLER_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16677_ _09156_ _09182_ _09319_ vssd1 vssd1 vccd1 vccd1 _09320_ sky130_fd_sc_hd__a21oi_1
X_13889_ _06621_ _06625_ _06576_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__o21a_1
XFILLER_59_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18416_ _01922_ _02114_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15628_ _05364_ _05461_ _07893_ vssd1 vssd1 vccd1 vccd1 _08273_ sky130_fd_sc_hd__mux2_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19396_ _02878_ _02881_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__xnor2_1
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18347_ _08802_ _01524_ _10139_ _09668_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__o22a_1
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15559_ _08202_ _08203_ vssd1 vssd1 vccd1 vccd1 _08204_ sky130_fd_sc_hd__and2_2
XFILLER_202_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18278_ _01870_ _01872_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__nor2_1
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput40 i_mode[2] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_4
X_17229_ _09804_ _09805_ _09806_ _09807_ vssd1 vssd1 vccd1 vccd1 _09808_ sky130_fd_sc_hd__a211o_1
XFILLER_190_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 i_vec_mosi vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_6
XFILLER_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21625_ clknet_leaf_28_i_clk _01394_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21556_ net477 _01325_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20507_ _03401_ _03402_ _03403_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__a21o_1
XFILLER_166_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21487_ net408 _01256_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_153_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11240_ gpout0.hpos\[3\] _04023_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__and2_1
XFILLER_5_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20438_ _03343_ _03344_ _03345_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__o21ai_1
XFILLER_175_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11171_ rbzero.otherx\[2\] _03929_ rbzero.map_rom.a6 _03958_ _03959_ vssd1 vssd1
+ vccd1 vccd1 _03960_ sky130_fd_sc_hd__o221a_1
XFILLER_101_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14930_ _07621_ _07628_ _07629_ _07620_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__o211a_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14861_ _05902_ _07426_ _07394_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__o21ai_1
XFILLER_169_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16600_ _08075_ vssd1 vssd1 vccd1 vccd1 _09243_ sky130_fd_sc_hd__buf_2
XFILLER_29_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13812_ _06426_ _06496_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__nor2_1
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17580_ _10124_ _10145_ vssd1 vssd1 vccd1 vccd1 _10146_ sky130_fd_sc_hd__xnor2_2
XFILLER_90_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14792_ _07487_ _07456_ _07522_ _07523_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__a211oi_4
XFILLER_204_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16531_ _09167_ _09174_ vssd1 vssd1 vccd1 vccd1 _09175_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13743_ _06475_ _06476_ _06477_ _06479_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__a22o_1
X_10955_ rbzero.tex_b1\[14\] rbzero.tex_b1\[15\] _03817_ vssd1 vssd1 vccd1 vccd1 _03825_
+ sky130_fd_sc_hd__mux2_1
XFILLER_113_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19250_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_sky\[3\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__mux2_1
XFILLER_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16462_ _09102_ _09105_ vssd1 vssd1 vccd1 vccd1 _09106_ sky130_fd_sc_hd__nor2_1
XFILLER_44_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ _06400_ _06404_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__nor2_1
X_10886_ rbzero.tex_b1\[47\] rbzero.tex_b1\[48\] _03784_ vssd1 vssd1 vccd1 vccd1 _03789_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18201_ _01802_ _01803_ _01901_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a21o_1
XFILLER_188_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15413_ _05209_ _08057_ vssd1 vssd1 vccd1 vccd1 _08058_ sky130_fd_sc_hd__or2_2
XFILLER_189_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12625_ rbzero.debug_overlay.playerY\[1\] _05378_ _05204_ vssd1 vssd1 vccd1 vccd1
+ _05379_ sky130_fd_sc_hd__mux2_1
X_19181_ rbzero.floor_leak\[1\] _02732_ _02735_ _02722_ vssd1 vssd1 vccd1 vccd1 _00741_
+ sky130_fd_sc_hd__o211a_1
X_16393_ _08352_ _08355_ _09036_ vssd1 vssd1 vccd1 vccd1 _09038_ sky130_fd_sc_hd__and3_1
XFILLER_106_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18132_ _01831_ _01832_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__or2_1
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15344_ _07988_ vssd1 vssd1 vccd1 vccd1 _07989_ sky130_fd_sc_hd__clkbuf_4
X_12556_ _05301_ _05305_ _05309_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__o21a_1
XFILLER_200_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11507_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _04273_ vssd1 vssd1 vccd1 vccd1 _04287_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18063_ _01762_ _01763_ _01755_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__a21o_1
XFILLER_145_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15275_ _07903_ _07918_ _07919_ vssd1 vssd1 vccd1 vccd1 _07920_ sky130_fd_sc_hd__a21o_1
X_12487_ rbzero.wall_tracer.trackDistX\[-11\] vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__inv_2
XFILLER_171_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17014_ _09618_ _09619_ _09653_ vssd1 vssd1 vccd1 vccd1 _09654_ sky130_fd_sc_hd__a21o_1
X_11438_ _04217_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__buf_6
X_14226_ _06805_ _06672_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__nor2_1
XFILLER_160_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14157_ _06805_ _06663_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__nor2_1
X_11369_ _04147_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__nand2_1
XFILLER_99_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13108_ _05814_ _05840_ _05843_ _05844_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__a22o_1
X_14088_ _06669_ _06824_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__xnor2_1
X_18965_ _02612_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__clkbuf_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17916_ _01498_ _08057_ _01618_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__or3_1
XFILLER_26_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _05759_ _05772_ _05775_ _05699_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__or4b_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18896_ rbzero.spi_registers.spi_counter\[2\] _02565_ vssd1 vssd1 vccd1 vccd1 _02566_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17847_ _10292_ _10295_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__nor2_1
XFILLER_120_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20208__231 clknet_1_0__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__inv_2
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17778_ _01473_ _01481_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__and2_1
XFILLER_82_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19517_ _02980_ _02994_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__nand2_1
X_16729_ _09364_ _09370_ vssd1 vssd1 vccd1 vccd1 _09371_ sky130_fd_sc_hd__xnor2_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19448_ _02913_ _02916_ _02929_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__and3_1
XFILLER_168_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19379_ _04034_ _02864_ _02865_ _02866_ _07706_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a221o_1
XFILLER_176_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21410_ net331 _01179_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21341_ net262 _01110_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20254__273 clknet_1_0__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__inv_2
XFILLER_118_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21272_ clknet_leaf_5_i_clk _01041_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_191_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20987_ clknet_leaf_12_i_clk _00756_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10740_ rbzero.tex_g0\[53\] rbzero.tex_g0\[52\] _03706_ vssd1 vssd1 vccd1 vccd1 _03712_
+ sky130_fd_sc_hd__mux2_1
XFILLER_81_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ rbzero.tex_g1\[21\] rbzero.tex_g1\[22\] _03669_ vssd1 vssd1 vccd1 vccd1 _03676_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ net36 _05165_ _05176_ net37 vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__o211a_1
XFILLER_22_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21608_ net149 _01377_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13390_ _06124_ _06125_ _06121_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__a21oi_1
XFILLER_90_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20337__348 clknet_1_0__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__inv_2
X_12341_ _05100_ _05106_ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__o21ai_1
XFILLER_167_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21539_ net460 _01308_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15060_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__nand2_1
X_12272_ _05035_ _05040_ net25 vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__and3b_1
XFILLER_175_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14011_ _06746_ _06747_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__nand2_1
X_11223_ _04007_ _04008_ _04009_ _03477_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__or4b_1
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03037_ clknet_0__03037_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03037_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_122_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ rbzero.debug_overlay.playerY\[1\] _03942_ vssd1 vssd1 vccd1 vccd1 _03943_
+ sky130_fd_sc_hd__nand2_1
XFILLER_175_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18750_ _02435_ _02436_ _02437_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__o21a_1
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11085_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _03887_ vssd1 vssd1 vccd1 vccd1 _03893_
+ sky130_fd_sc_hd__mux2_1
X_15962_ _08587_ _08604_ vssd1 vssd1 vccd1 vccd1 _08607_ sky130_fd_sc_hd__nor2_1
XFILLER_23_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17701_ _10139_ vssd1 vssd1 vccd1 vccd1 _10266_ sky130_fd_sc_hd__clkbuf_4
X_14913_ rbzero.wall_tracer.trackDistY\[-3\] rbzero.wall_tracer.trackDistX\[-3\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__mux2_1
X_18681_ _02293_ _02298_ _02376_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a21o_1
XFILLER_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _08535_ _08536_ _08537_ vssd1 vssd1 vccd1 vccd1 _08538_ sky130_fd_sc_hd__a21oi_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ _10069_ _10083_ _10196_ vssd1 vssd1 vccd1 vccd1 _10197_ sky130_fd_sc_hd__a21o_1
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14844_ _07565_ vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__clkbuf_1
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20082__118 clknet_1_0__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__inv_2
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17563_ _05211_ _09699_ _10128_ vssd1 vssd1 vccd1 vccd1 _10129_ sky130_fd_sc_hd__o21a_1
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14775_ _07477_ _07479_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__nor2_1
XFILLER_95_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11987_ _04247_ _04759_ _04760_ _04761_ _04254_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__o221a_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19302_ rbzero.spi_registers.new_other\[6\] rbzero.spi_registers.spi_buffer\[6\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__mux2_1
X_16514_ _09040_ _08430_ _09041_ _09157_ vssd1 vssd1 vccd1 vccd1 _09158_ sky130_fd_sc_hd__o31ai_4
X_13726_ _06426_ _06462_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__nor2_1
XFILLER_32_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17494_ _10058_ _10059_ vssd1 vssd1 vccd1 vccd1 _10060_ sky130_fd_sc_hd__nand2_1
X_10938_ rbzero.tex_b1\[22\] rbzero.tex_b1\[23\] _03806_ vssd1 vssd1 vccd1 vccd1 _03816_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19233_ rbzero.spi_registers.new_vshift\[3\] _02763_ vssd1 vssd1 vccd1 vccd1 _02768_
+ sky130_fd_sc_hd__or2_1
XFILLER_108_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16445_ _09056_ _09058_ vssd1 vssd1 vccd1 vccd1 _09089_ sky130_fd_sc_hd__nand2_1
X_10869_ rbzero.tex_b1\[55\] rbzero.tex_b1\[56\] _03773_ vssd1 vssd1 vccd1 vccd1 _03780_
+ sky130_fd_sc_hd__mux2_1
X_13657_ _06388_ _06390_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19164_ rbzero.othery\[2\] _02710_ _02723_ _02722_ vssd1 vssd1 vccd1 vccd1 _00736_
+ sky130_fd_sc_hd__o211a_1
X_12608_ _05308_ _05312_ _05318_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__o21ai_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _09000_ _09020_ vssd1 vssd1 vccd1 vccd1 _09021_ sky130_fd_sc_hd__xnor2_4
X_13588_ _06281_ _06283_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__nor2_1
X_18115_ _01814_ _01815_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__nor2_1
XFILLER_9_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15327_ _07971_ _05488_ vssd1 vssd1 vccd1 vccd1 _07972_ sky130_fd_sc_hd__nor2_1
XFILLER_173_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19095_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.spi_buffer\[2\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__mux2_1
X_12539_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] _05291_
+ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__a31o_1
XFILLER_185_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18046_ _01746_ _01747_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__xor2_1
XFILLER_133_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15258_ rbzero.wall_tracer.state\[13\] vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__clkbuf_4
XFILLER_144_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14209_ _06932_ _06945_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__or2b_1
X_15189_ rbzero.wall_tracer.rayAddendX\[6\] rbzero.wall_tracer.rayAddendX\[5\] rbzero.wall_tracer.rayAddendX\[4\]
+ rbzero.wall_tracer.rayAddendX\[3\] _07785_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__o41a_1
XFILLER_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19997_ rbzero.pov.ready_buffer\[1\] _03239_ _03242_ rbzero.debug_overlay.vplaneY\[-8\]
+ _03254_ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__o221a_1
XFILLER_154_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18948_ _02603_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18879_ rbzero.wall_tracer.trackDistY\[11\] rbzero.wall_tracer.stepDistY\[11\] vssd1
+ vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__xor2_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20910_ clknet_leaf_78_i_clk _00679_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_20284__299 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__inv_2
XFILLER_54_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20841_ clknet_leaf_62_i_clk _00610_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20772_ clknet_leaf_40_i_clk _00541_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21324_ net245 _01093_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_198_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21255_ clknet_leaf_84_i_clk _01024_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_144_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21186_ clknet_leaf_74_i_clk _00955_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11910_ _04684_ _04685_ _04265_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__mux2_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _05562_ _05565_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__and2_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _04230_ _04613_ _04617_ _04232_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a211o_1
XFILLER_166_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _04129_ vssd1 vssd1 vccd1 vccd1 _04550_
+ sky130_fd_sc_hd__mux2_1
X_14560_ _07291_ _07296_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__nand2_1
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10723_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _03624_ vssd1 vssd1 vccd1 vccd1 _03703_
+ sky130_fd_sc_hd__mux2_1
X_13511_ _06237_ _06238_ _06247_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__a21oi_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14491_ _07137_ _07045_ _07166_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__a21o_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _08871_ _08874_ vssd1 vssd1 vccd1 vccd1 _08875_ sky130_fd_sc_hd__nor2_1
X_10654_ rbzero.tex_g1\[29\] rbzero.tex_g1\[30\] _03658_ vssd1 vssd1 vccd1 vccd1 _03667_
+ sky130_fd_sc_hd__mux2_1
X_13442_ _06078_ _06067_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__or2_1
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13373_ _06037_ _06092_ _06108_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__a21oi_1
X_16161_ _08737_ _08761_ vssd1 vssd1 vccd1 vccd1 _08806_ sky130_fd_sc_hd__xnor2_2
X_10585_ _03630_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15112_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__or2_1
X_12324_ _05087_ _04738_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__nor2_1
X_16092_ _08725_ _08734_ _08736_ vssd1 vssd1 vccd1 vccd1 _08737_ sky130_fd_sc_hd__a21oi_2
XFILLER_86_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12255_ net23 net24 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__nand2_1
XFILLER_181_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15043_ _07703_ _07704_ _07705_ _07706_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__a31o_1
X_19920_ _03216_ _03217_ _02822_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__a21oi_1
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11206_ _03933_ rbzero.map_rom.i_row\[4\] _03990_ _03994_ vssd1 vssd1 vccd1 vccd1
+ _03995_ sky130_fd_sc_hd__or4_1
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19851_ rbzero.pov.ready_buffer\[67\] _03164_ vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__nor2_1
X_12186_ _04904_ _04925_ _04956_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__a21oi_2
XFILLER_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11137_ rbzero.debug_overlay.playerX\[1\] vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__inv_2
X_18802_ _05532_ _02483_ _02484_ _02399_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__o31a_1
XFILLER_205_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19782_ rbzero.pov.spi_buffer\[64\] rbzero.pov.spi_buffer\[65\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03120_ sky130_fd_sc_hd__mux2_1
X_16994_ _09631_ _09632_ vssd1 vssd1 vccd1 vccd1 _09634_ sky130_fd_sc_hd__nand2_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18733_ _02421_ _02422_ _02423_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__nor3_1
X_11068_ rbzero.tex_b0\[25\] rbzero.tex_b0\[24\] _03876_ vssd1 vssd1 vccd1 vccd1 _03884_
+ sky130_fd_sc_hd__mux2_1
X_15945_ _08522_ _08523_ vssd1 vssd1 vccd1 vccd1 _08590_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18664_ _08257_ _09215_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__nor2_1
XFILLER_110_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15876_ _07601_ _04014_ _05197_ _07992_ vssd1 vssd1 vccd1 vccd1 _08521_ sky130_fd_sc_hd__and4_1
XFILLER_110_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17615_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] vssd1
+ vssd1 vccd1 vccd1 _10180_ sky130_fd_sc_hd__nor2_1
X_14827_ rbzero.wall_tracer.stepDistY\[-1\] _07461_ vssd1 vssd1 vccd1 vccd1 _07553_
+ sky130_fd_sc_hd__nor2_1
X_18595_ _02198_ _02164_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__or2b_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17546_ _09686_ _09980_ _10111_ vssd1 vssd1 vccd1 vccd1 _10112_ sky130_fd_sc_hd__a21bo_1
XFILLER_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14758_ _07477_ _07489_ _07491_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__a21oi_1
XFILLER_205_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13709_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__or2_1
XFILLER_60_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17477_ _09933_ _09936_ _10041_ vssd1 vssd1 vccd1 vccd1 _10043_ sky130_fd_sc_hd__and3_1
X_14689_ _07106_ _07425_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__or2_1
XFILLER_177_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19216_ rbzero.spi_registers.new_floor\[3\] rbzero.spi_registers.got_new_floor _02711_
+ _03911_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a31o_1
X_16428_ _09071_ _09069_ _09070_ vssd1 vssd1 vccd1 vccd1 _09073_ sky130_fd_sc_hd__and3_1
XFILLER_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19147_ _05190_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__clkbuf_4
XFILLER_146_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16359_ _07967_ _08035_ _08046_ _08674_ vssd1 vssd1 vccd1 vccd1 _09004_ sky130_fd_sc_hd__o22ai_1
XFILLER_9_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19078_ _02671_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18029_ _01715_ _01730_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__xnor2_1
XFILLER_160_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21040_ clknet_leaf_77_i_clk _00809_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20366__374 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__inv_2
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20065__102 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__inv_2
XFILLER_55_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20824_ clknet_leaf_48_i_clk _00593_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20755_ clknet_leaf_40_i_clk _00524_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20686_ clknet_leaf_64_i_clk _00470_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ _03515_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21307_ net228 _01076_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_105_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _04163_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__clkbuf_4
X_21238_ clknet_leaf_79_i_clk _01007_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19609__63 clknet_1_1__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__inv_2
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21169_ clknet_leaf_92_i_clk _00938_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19624__77 clknet_1_0__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__inv_2
XFILLER_65_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13991_ _06698_ _06726_ _06671_ _06727_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__o31a_1
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _08302_ _08374_ vssd1 vssd1 vccd1 vccd1 _08375_ sky130_fd_sc_hd__xor2_1
XFILLER_86_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _05604_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__clkinv_2
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _08299_ _08305_ vssd1 vssd1 vccd1 vccd1 _08306_ sky130_fd_sc_hd__xor2_1
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _04000_ _05488_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nand2_1
XFILLER_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17400_ _09965_ _09966_ vssd1 vssd1 vccd1 vccd1 _09967_ sky130_fd_sc_hd__xnor2_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _07218_ _07323_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__xor2_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18380_ _02075_ _02077_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__nand2_1
X_11824_ _04597_ _04600_ _04332_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__mux2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _08231_ _08236_ _05209_ vssd1 vssd1 vccd1 vccd1 _08237_ sky130_fd_sc_hd__a21o_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _09899_ sky130_fd_sc_hd__and2_1
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _07160_ _07199_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__xor2_1
XFILLER_53_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _04531_ _04532_ _04138_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__mux2_1
XFILLER_202_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10706_ _03694_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17262_ _09837_ vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14474_ _07203_ _07210_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11686_ _04430_ _04431_ _04450_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__and3_2
XFILLER_144_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19001_ _02631_ vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16213_ _08855_ _08857_ vssd1 vssd1 vccd1 vccd1 _08858_ sky130_fd_sc_hd__nand2_1
XFILLER_128_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13425_ _05978_ _06161_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__nor2_1
X_10637_ _03646_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__clkbuf_4
X_17193_ _09774_ _09776_ vssd1 vssd1 vccd1 vccd1 _09778_ sky130_fd_sc_hd__nand2_1
X_16144_ _08769_ _08788_ vssd1 vssd1 vccd1 vccd1 _08789_ sky130_fd_sc_hd__xnor2_1
X_10568_ _03621_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13356_ _05945_ _05949_ _05939_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__a21oi_1
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12307_ _05062_ _05075_ _05035_ net25 vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__o211a_1
XFILLER_143_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16075_ _07989_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08720_ sky130_fd_sc_hd__or3_2
XFILLER_127_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10499_ _03585_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__clkbuf_1
X_13287_ _06010_ _06012_ _06023_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__a21o_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15026_ _07684_ _07689_ _07690_ vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__o21ai_2
X_19903_ rbzero.pov.ready_buffer\[48\] _02823_ _03193_ _03205_ vssd1 vssd1 vccd1 vccd1
+ _03206_ sky130_fd_sc_hd__a211o_1
X_12238_ _04996_ _05005_ _04986_ _05007_ net19 vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__o2111a_1
XFILLER_155_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ _04907_ _04905_ _04938_ _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__a31o_1
X_19834_ _07901_ _03143_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__nand2_1
XFILLER_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16977_ _09498_ _09512_ _09510_ vssd1 vssd1 vccd1 vccd1 _09617_ sky130_fd_sc_hd__a21o_1
X_19765_ rbzero.pov.spi_buffer\[56\] rbzero.pov.spi_buffer\[57\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03111_ sky130_fd_sc_hd__mux2_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput5 i_gpout0_sel[3] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_8
XFILLER_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15928_ _08096_ _08572_ vssd1 vssd1 vccd1 vccd1 _08573_ sky130_fd_sc_hd__or2_1
X_18716_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__and2_1
X_19696_ rbzero.pov.spi_buffer\[23\] rbzero.pov.spi_buffer\[24\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03075_ sky130_fd_sc_hd__mux2_1
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18647_ _10248_ _02150_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__and2_1
Xclkbuf_0__03296_ _03296_ vssd1 vssd1 vccd1 vccd1 clknet_0__03296_ sky130_fd_sc_hd__clkbuf_16
X_15859_ _08496_ _08502_ vssd1 vssd1 vccd1 vccd1 _08504_ sky130_fd_sc_hd__nor2_1
XFILLER_65_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18578_ _02273_ _02274_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__xor2_1
XFILLER_206_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17529_ _08178_ _08493_ _08044_ _10094_ vssd1 vssd1 vccd1 vccd1 _10095_ sky130_fd_sc_hd__o22ai_1
XFILLER_33_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20540_ rbzero.traced_texa\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03431_
+ sky130_fd_sc_hd__nand2_1
XFILLER_123_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20471_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 _03373_
+ sky130_fd_sc_hd__and2_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21023_ clknet_leaf_3_i_clk _00792_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20807_ clknet_leaf_25_i_clk _00576_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ gpout0.vpos\[2\] gpout0.vpos\[1\] gpout0.vpos\[0\] _04319_ vssd1 vssd1 vccd1
+ vccd1 _04320_ sky130_fd_sc_hd__o31a_4
X_20738_ clknet_3_5_0_i_clk _00507_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11471_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _04250_ vssd1 vssd1 vccd1 vccd1 _04251_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20669_ clknet_leaf_61_i_clk _00453_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10422_ rbzero.tex_r1\[9\] rbzero.tex_r1\[10\] _03538_ vssd1 vssd1 vccd1 vccd1 _03543_
+ sky130_fd_sc_hd__mux2_1
X_13210_ _05865_ _05870_ _05875_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nor3b_1
XFILLER_109_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14190_ _06769_ _06677_ _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__o21ba_1
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10353_ rbzero.tex_r1\[42\] rbzero.tex_r1\[43\] _03505_ vssd1 vssd1 vccd1 vccd1 _03507_
+ sky130_fd_sc_hd__mux2_1
X_13141_ _05827_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__clkinv_2
XFILLER_136_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ _05740_ _05777_ _05790_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__or3_1
XFILLER_183_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16900_ _08170_ _09419_ _09540_ vssd1 vssd1 vccd1 vccd1 _09541_ sky130_fd_sc_hd__or3_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12023_ rbzero.tex_b1\[35\] rbzero.tex_b1\[34\] _04337_ vssd1 vssd1 vccd1 vccd1 _04798_
+ sky130_fd_sc_hd__mux2_1
X_17880_ _09522_ _09029_ _01582_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__or3_1
XFILLER_151_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16831_ _09352_ _09361_ vssd1 vssd1 vccd1 vccd1 _09472_ sky130_fd_sc_hd__or2b_1
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19550_ rbzero.pov.spi_counter\[0\] _03019_ rbzero.pov.spi_counter\[1\] vssd1 vssd1
+ vccd1 vccd1 _03023_ sky130_fd_sc_hd__a21o_1
X_16762_ _09386_ _09403_ vssd1 vssd1 vccd1 vccd1 _09404_ sky130_fd_sc_hd__xor2_1
XFILLER_150_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13974_ _06031_ _06707_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__nor2_1
XFILLER_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18501_ _02164_ _02198_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15713_ _08355_ _08357_ vssd1 vssd1 vccd1 vccd1 _08358_ sky130_fd_sc_hd__and2_1
X_19481_ _02905_ rbzero.debug_overlay.vplaneY\[-2\] vssd1 vssd1 vccd1 vccd1 _02961_
+ sky130_fd_sc_hd__nor2_1
X_12925_ _05650_ _05655_ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__or3_1
XFILLER_207_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16693_ _09334_ _09335_ vssd1 vssd1 vccd1 vccd1 _09336_ sky130_fd_sc_hd__or2b_1
XFILLER_111_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18432_ _02128_ _02130_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__nand2_1
XFILLER_62_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15644_ _08191_ _08265_ _08277_ _08267_ vssd1 vssd1 vccd1 vccd1 _08289_ sky130_fd_sc_hd__a22o_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12856_ rbzero.wall_tracer.rayAddendX\[-3\] _05592_ _05560_ vssd1 vssd1 vccd1 vccd1
+ _05593_ sky130_fd_sc_hd__mux2_2
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _01951_ _01963_ _02061_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__a21o_1
X_20202__226 clknet_1_1__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__inv_2
X_11807_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _04341_ vssd1 vssd1 vccd1 vccd1 _04585_
+ sky130_fd_sc_hd__mux2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15575_ _07560_ _07562_ _07564_ _08171_ vssd1 vssd1 vccd1 vccd1 _08220_ sky130_fd_sc_hd__or4_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _05530_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_199_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _09880_ _09881_ _09882_ vssd1 vssd1 vccd1 vccd1 _09884_ sky130_fd_sc_hd__a21oi_1
XFILLER_187_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14526_ _07070_ _07079_ _07262_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__a21oi_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18294_ _01992_ _01993_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__xor2_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11738_ _04510_ _04516_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__or2_1
XFILLER_159_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17245_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _09822_ sky130_fd_sc_hd__nand2_1
X_14457_ _07184_ _07193_ _07191_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11669_ _04422_ _04447_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__nand2_2
X_13408_ _06091_ _06144_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__and2b_1
XFILLER_179_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17176_ rbzero.traced_texa\[4\] _09770_ _09769_ rbzero.wall_tracer.visualWallDist\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__a22o_1
X_14388_ _07122_ _07124_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__or2b_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16127_ _08768_ _08770_ _08771_ vssd1 vssd1 vccd1 vccd1 _08772_ sky130_fd_sc_hd__o21a_1
XFILLER_128_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13339_ _06044_ _06047_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__and2b_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16058_ _07601_ _08148_ _07990_ _07962_ vssd1 vssd1 vccd1 vccd1 _08703_ sky130_fd_sc_hd__and4_1
XFILLER_130_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15009_ rbzero.wall_tracer.stepDistX\[11\] _07589_ _05201_ vssd1 vssd1 vccd1 vccd1
+ _07675_ sky130_fd_sc_hd__mux2_1
XFILLER_130_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19817_ _03138_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__clkbuf_4
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03317_ clknet_0__03317_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03317_
+ sky130_fd_sc_hd__clkbuf_16
X_19748_ rbzero.pov.spi_buffer\[48\] rbzero.pov.spi_buffer\[49\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03102_ sky130_fd_sc_hd__mux2_1
X_19603__58 clknet_1_1__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__inv_2
XFILLER_37_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19679_ rbzero.pov.spi_buffer\[15\] rbzero.pov.spi_buffer\[16\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03066_ sky130_fd_sc_hd__mux2_1
XFILLER_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21641_ clknet_leaf_29_i_clk _01410_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20177__203 clknet_1_0__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__inv_2
Xclkbuf_opt_6_0_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_6_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_162_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21572_ net493 _01341_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[23\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_10 _07541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_21 _09765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20523_ rbzero.traced_texa\[6\] rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _03417_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_43 _07536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_65 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_76 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20454_ _03351_ _03355_ _03352_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__o21ai_1
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_84_i_clk clknet_opt_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21006_ clknet_leaf_9_i_clk _00775_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_101_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ _03833_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12710_ _05416_ _05442_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__nand2_1
X_13690_ _06394_ _06416_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_22_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_188_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12641_ _05391_ _05392_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15360_ _08004_ rbzero.debug_overlay.playerY\[-7\] _05374_ vssd1 vssd1 vccd1 vccd1
+ _08005_ sky130_fd_sc_hd__mux2_2
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[11\] vssd1
+ vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__nand2_1
XFILLER_106_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14311_ _06067_ _06678_ _07047_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__or3b_1
X_11523_ rbzero.tex_r0\[31\] _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__and3_1
XFILLER_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_i_clk clknet_opt_8_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15291_ _07933_ _07536_ _07935_ vssd1 vssd1 vccd1 vccd1 _07936_ sky130_fd_sc_hd__o21ai_4
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17030_ _09276_ _08111_ vssd1 vssd1 vccd1 vccd1 _09670_ sky130_fd_sc_hd__nor2_4
XFILLER_172_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14242_ _06967_ _06968_ _06976_ _06978_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__a211oi_1
X_11454_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _04214_ vssd1 vssd1 vccd1 vccd1 _04234_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10405_ rbzero.tex_r1\[17\] rbzero.tex_r1\[18\] _03527_ vssd1 vssd1 vccd1 vccd1 _03534_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11385_ rbzero.row_render.size\[0\] vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__inv_2
X_14173_ _06887_ _06901_ _06909_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__o21a_1
XFILLER_152_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13124_ _05645_ _05796_ _05860_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__o21ai_1
XFILLER_113_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10336_ rbzero.tex_r1\[50\] rbzero.tex_r1\[51\] _03494_ vssd1 vssd1 vccd1 vccd1 _03498_
+ sky130_fd_sc_hd__mux2_1
X_18981_ rbzero.pov.spi_buffer\[23\] rbzero.pov.ready_buffer\[23\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02621_ sky130_fd_sc_hd__mux2_1
XFILLER_112_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17932_ _10134_ _10131_ _01527_ _01525_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__a31o_1
XFILLER_124_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _05791_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12006_ _04779_ _04780_ _04304_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__mux2_1
X_17863_ _01563_ _01565_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__nand2_1
XFILLER_39_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16814_ _09454_ _09455_ vssd1 vssd1 vccd1 vccd1 _09456_ sky130_fd_sc_hd__or2_2
XFILLER_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xnet99_4 clknet_1_1__leaf__04835_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__inv_2
X_17794_ _08188_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__clkbuf_4
XFILLER_207_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16745_ _07996_ _08705_ _08035_ _08046_ vssd1 vssd1 vccd1 vccd1 _09387_ sky130_fd_sc_hd__or4_1
X_19533_ _02906_ _04034_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__or3_1
X_13957_ _06681_ _06688_ _06691_ _06693_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19464_ _02944_ _02945_ _04029_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__o21ai_1
X_12908_ _05618_ _05644_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__xor2_2
XFILLER_207_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16676_ _09153_ _09155_ vssd1 vssd1 vccd1 vccd1 _09319_ sky130_fd_sc_hd__nor2_1
XFILLER_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13888_ _06622_ _06624_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18415_ _02112_ _02113_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__and2_1
XFILLER_185_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15627_ _07549_ _08270_ _08271_ _07933_ vssd1 vssd1 vccd1 vccd1 _08272_ sky130_fd_sc_hd__a211o_2
XFILLER_22_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19395_ _02879_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__nand2_1
XFILLER_72_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ rbzero.wall_tracer.visualWallDist\[10\] _05571_ _05572_ vssd1 vssd1 vccd1
+ vccd1 _05576_ sky130_fd_sc_hd__a21o_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18346_ _08802_ _09668_ _01524_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__or3_2
XFILLER_194_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15558_ _05208_ rbzero.wall_tracer.stepDistX\[0\] vssd1 vssd1 vccd1 vccd1 _08203_
+ sky130_fd_sc_hd__nand2_2
XFILLER_33_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14509_ _07235_ _07244_ _07245_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__a21oi_1
X_18277_ _01975_ _01976_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__nor2_1
XFILLER_175_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15489_ _04013_ rbzero.wall_tracer.stepDistY\[-12\] vssd1 vssd1 vccd1 vccd1 _08134_
+ sky130_fd_sc_hd__or2_1
XFILLER_200_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17228_ _05203_ vssd1 vssd1 vccd1 vccd1 _09807_ sky130_fd_sc_hd__buf_6
XFILLER_163_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput30 i_gpout4_sel[4] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_6
XFILLER_174_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput41 i_reg_csb vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_16
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput52 i_vec_sclk vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_8
XFILLER_162_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17159_ rbzero.traced_texa\[-10\] _09766_ _09767_ _07601_ vssd1 vssd1 vccd1 vccd1
+ _00547_ sky130_fd_sc_hd__a22o_1
XFILLER_115_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21624_ clknet_leaf_27_i_clk _01393_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_179_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21555_ net476 _01324_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20506_ _03396_ _03399_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__nand2_1
X_21486_ net407 _01255_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20437_ _03338_ _03341_ _03339_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__a21boi_1
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11170_ rbzero.otherx\[2\] _03929_ _03935_ rbzero.othery\[4\] vssd1 vssd1 vccd1 vccd1
+ _03959_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20231__252 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__inv_2
XFILLER_136_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14860_ _07433_ _07445_ _07446_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__nor3_1
XFILLER_169_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13811_ _06497_ _06498_ _06547_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14791_ _07511_ _07437_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__nor2_1
XFILLER_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ _09168_ _09173_ vssd1 vssd1 vccd1 vccd1 _09174_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13742_ _06475_ _06478_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__xnor2_1
X_19594__49 clknet_1_1__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__inv_2
XFILLER_204_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10954_ _03824_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16461_ _07941_ _09103_ _09010_ _09104_ vssd1 vssd1 vccd1 vccd1 _09105_ sky130_fd_sc_hd__o31a_1
XFILLER_204_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13673_ _06408_ _06409_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__xor2_1
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10885_ _03788_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__clkbuf_1
X_18200_ _01804_ _01900_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__xor2_1
XFILLER_189_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15412_ rbzero.wall_tracer.visualWallDist\[2\] _04015_ vssd1 vssd1 vccd1 vccd1 _08057_
+ sky130_fd_sc_hd__nand2_2
XFILLER_176_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12624_ _03925_ _05377_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__xnor2_1
X_19180_ rbzero.spi_registers.new_leak\[1\] _02733_ vssd1 vssd1 vccd1 vccd1 _02735_
+ sky130_fd_sc_hd__or2_1
X_16392_ _08352_ _08355_ _09036_ vssd1 vssd1 vccd1 vccd1 _09037_ sky130_fd_sc_hd__a21oi_1
XFILLER_169_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18131_ _01582_ _01706_ _01708_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__o21a_1
XFILLER_129_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15343_ _05206_ _07984_ _07987_ vssd1 vssd1 vccd1 vccd1 _07988_ sky130_fd_sc_hd__o21ai_4
X_12555_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__or2_1
XFILLER_196_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18062_ _01755_ _01762_ _01763_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__nand3_1
X_11506_ rbzero.tex_r0\[2\] _04214_ _04219_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__a21o_1
X_15274_ rbzero.wall_tracer.visualWallDist\[-5\] _04012_ rbzero.wall_tracer.state\[6\]
+ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__a21o_1
XFILLER_157_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ rbzero.wall_tracer.trackDistX\[-10\] vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__inv_2
XFILLER_144_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17013_ _09638_ _09652_ vssd1 vssd1 vccd1 vccd1 _09653_ sky130_fd_sc_hd__xnor2_1
X_20314__327 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__inv_2
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14225_ _06946_ _06949_ _06961_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__a21oi_1
X_11437_ _04125_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__buf_6
XFILLER_99_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14156_ _06865_ _06867_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__xnor2_1
X_11368_ rbzero.row_render.size\[1\] rbzero.row_render.size\[0\] vssd1 vssd1 vccd1
+ vccd1 _04148_ sky130_fd_sc_hd__nor2_1
XFILLER_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13107_ _05811_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__clkbuf_4
XFILLER_112_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10319_ rbzero.tex_r1\[58\] rbzero.tex_r1\[59\] _03483_ vssd1 vssd1 vccd1 vccd1 _03489_
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14087_ _06666_ _06668_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__nor2_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ rbzero.pov.spi_buffer\[15\] rbzero.pov.ready_buffer\[15\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02612_ sky130_fd_sc_hd__mux2_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11299_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] vssd1 vssd1
+ vccd1 vccd1 _04079_ sky130_fd_sc_hd__nand2_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _01616_ _01617_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _05684_ _05689_ _05703_ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18895_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\] _02564_
+ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__a21o_1
XFILLER_152_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17846_ _01548_ _01549_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__nor2_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17777_ _01479_ _01480_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14989_ rbzero.wall_tracer.stepDistX\[1\] _07560_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07665_ sky130_fd_sc_hd__mux2_1
XFILLER_75_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19516_ _02905_ rbzero.debug_overlay.vplaneY\[0\] vssd1 vssd1 vccd1 vccd1 _02994_
+ sky130_fd_sc_hd__or2_1
X_16728_ _09367_ _09369_ vssd1 vssd1 vccd1 vccd1 _09370_ sky130_fd_sc_hd__xor2_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16659_ _09132_ _09144_ _09301_ vssd1 vssd1 vccd1 vccd1 _09302_ sky130_fd_sc_hd__a21bo_1
X_19447_ _02913_ _02916_ _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19378_ rbzero.debug_overlay.vplaneY\[-6\] _02849_ _04034_ vssd1 vssd1 vccd1 vccd1
+ _02866_ sky130_fd_sc_hd__a21oi_1
XFILLER_33_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18329_ _01971_ _02027_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__xor2_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21340_ net261 _01109_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21271_ clknet_leaf_5_i_clk _01040_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
X_20289__304 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__inv_2
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20986_ clknet_leaf_9_i_clk _00755_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10670_ _03675_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21607_ net148 _01376_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12340_ net41 _05084_ _05107_ net43 net29 vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__a221o_1
XFILLER_139_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21538_ net459 _01307_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12271_ _05036_ _05037_ _05038_ _05039_ net22 net21 vssd1 vssd1 vccd1 vccd1 _05040_
+ sky130_fd_sc_hd__mux4_1
XFILLER_175_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21469_ net390 _01238_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14010_ _06680_ _06662_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__nor2_1
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11222_ gpout0.hpos\[7\] gpout0.hpos\[8\] vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__or2_1
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11153_ rbzero.map_rom.c6 vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__buf_2
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15961_ _08582_ _08568_ vssd1 vssd1 vccd1 vccd1 _08606_ sky130_fd_sc_hd__xnor2_2
X_11084_ _03892_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17700_ _09117_ _09991_ vssd1 vssd1 vccd1 vccd1 _10265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14912_ _05278_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__buf_4
XFILLER_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18680_ _02208_ _02299_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__and2b_1
X_15892_ _08513_ _08534_ vssd1 vssd1 vccd1 vccd1 _08537_ sky130_fd_sc_hd__nor2_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ _10080_ _10082_ vssd1 vssd1 vccd1 vccd1 _10196_ sky130_fd_sc_hd__nor2_1
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14843_ rbzero.wall_tracer.stepDistY\[3\] _07564_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07565_ sky130_fd_sc_hd__mux2_1
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17562_ _05211_ rbzero.wall_tracer.stepDistX\[11\] vssd1 vssd1 vccd1 vccd1 _10128_
+ sky130_fd_sc_hd__nand2_2
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14774_ _07477_ _07470_ _07506_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ rbzero.tex_b1\[10\] _04273_ _04304_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a21o_1
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16513_ _09030_ _09043_ vssd1 vssd1 vccd1 vccd1 _09157_ sky130_fd_sc_hd__nand2_1
XFILLER_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19301_ _02806_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13725_ _06458_ _06460_ _06461_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__a21o_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17493_ _09245_ _09243_ _09028_ _09164_ vssd1 vssd1 vccd1 vccd1 _10059_ sky130_fd_sc_hd__or4_1
X_10937_ _03815_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16444_ _08549_ _08957_ _09060_ _09087_ vssd1 vssd1 vccd1 vccd1 _09088_ sky130_fd_sc_hd__a31o_1
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19232_ rbzero.spi_registers.vshift\[2\] _02762_ _02767_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00760_ sky130_fd_sc_hd__o211a_1
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ _06350_ _06392_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__xnor2_1
XFILLER_182_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10868_ _03779_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ _05351_ _05353_ _05356_ _05360_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__or4_1
X_19163_ rbzero.spi_registers.new_other\[2\] _02712_ vssd1 vssd1 vccd1 vccd1 _02723_
+ sky130_fd_sc_hd__or2_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _09002_ _09019_ vssd1 vssd1 vccd1 vccd1 _09020_ sky130_fd_sc_hd__xnor2_2
XFILLER_129_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13587_ _06304_ _06323_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__nand2_1
XFILLER_185_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10799_ _03743_ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__clkbuf_1
X_18114_ _01805_ _01806_ _01813_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__and3_1
XFILLER_185_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15326_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__inv_2
XFILLER_184_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19094_ _02680_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__clkbuf_1
X_12538_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__and2_1
XFILLER_158_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18045_ _09674_ _09973_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__nor2_1
X_15257_ _07900_ _07901_ _05495_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__mux2_1
XFILLER_172_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12469_ rbzero.wall_tracer.trackDistX\[4\] vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__inv_2
XFILLER_160_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14208_ _06934_ _06939_ _06944_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__o21ai_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15188_ _07818_ _07819_ _07828_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__nor3_1
XFILLER_141_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14139_ _06859_ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19996_ rbzero.pov.ready_buffer\[0\] _03252_ _03253_ rbzero.debug_overlay.vplaneY\[-9\]
+ _03254_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__o221a_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18947_ rbzero.pov.spi_buffer\[7\] rbzero.pov.ready_buffer\[7\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02603_ sky130_fd_sc_hd__mux2_1
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18878_ _02546_ _02547_ _02545_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__o21ai_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17829_ _01530_ _01531_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__nand2_1
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20840_ clknet_leaf_58_i_clk _00609_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_165_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20771_ clknet_leaf_39_i_clk _00540_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21323_ net244 _01092_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21254_ clknet_leaf_87_i_clk _01023_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_2_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20205_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__buf_1
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21185_ clknet_leaf_74_i_clk _00954_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20343__353 clknet_1_0__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__inv_2
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _04379_ _04614_ _04615_ _04616_ _04209_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__o221a_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _04547_ _04548_ _04126_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__mux2_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20969_ clknet_leaf_7_i_clk _00738_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ _06244_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__nand2_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10722_ _03702_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14490_ _07220_ _07226_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__xor2_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ _06083_ _06086_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__and2b_1
X_10653_ _03666_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16160_ _08803_ _08804_ vssd1 vssd1 vccd1 vccd1 _08805_ sky130_fd_sc_hd__or2_1
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13372_ _06037_ _06092_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__and3_1
X_10584_ rbzero.tex_g1\[62\] rbzero.tex_g1\[63\] _03549_ vssd1 vssd1 vccd1 vccd1 _03630_
+ sky130_fd_sc_hd__mux2_1
XFILLER_194_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15111_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__nand2_1
X_12323_ net29 net30 vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__nand2_1
XFILLER_126_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16091_ _08661_ _08735_ vssd1 vssd1 vccd1 vccd1 _08736_ sky130_fd_sc_hd__or2_1
XFILLER_5_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15042_ _07695_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__buf_4
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12254_ _05021_ net61 _05022_ net24 vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__o211a_1
XFILLER_182_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11205_ rbzero.map_rom.f4 rbzero.map_rom.d6 _03921_ _03977_ vssd1 vssd1 vccd1 vccd1
+ _03994_ sky130_fd_sc_hd__or4_1
XFILLER_122_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19850_ _03146_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__clkbuf_4
X_12185_ _04930_ _04934_ _04942_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__o31a_1
X_18801_ _02480_ _02481_ _02479_ _02476_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__o211a_1
X_11136_ rbzero.map_rom.d6 vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__clkinv_2
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19781_ _03119_ vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16993_ _09631_ _09632_ vssd1 vssd1 vccd1 vccd1 _09633_ sky130_fd_sc_hd__or2_1
XFILLER_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18732_ _02414_ _02416_ _02415_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a21boi_1
X_11067_ _03883_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15944_ _08555_ _08554_ vssd1 vssd1 vccd1 vccd1 _08589_ sky130_fd_sc_hd__xor2_2
XFILLER_114_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18663_ _02354_ _02358_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__xnor2_1
X_15875_ _07974_ _08519_ vssd1 vssd1 vccd1 vccd1 _08520_ sky130_fd_sc_hd__nor2_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14826_ _07486_ _07455_ _07551_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__a21oi_4
XFILLER_97_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17614_ rbzero.wall_tracer.trackDistX\[2\] rbzero.wall_tracer.stepDistX\[2\] vssd1
+ vssd1 vccd1 vccd1 _10179_ sky130_fd_sc_hd__and2_1
XFILLER_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18594_ _02288_ _02290_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__xnor2_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ _10110_ _09417_ _09982_ vssd1 vssd1 vccd1 vccd1 _10111_ sky130_fd_sc_hd__or3_1
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14757_ _07477_ _07490_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__nor2_1
XFILLER_45_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11969_ _04742_ _04743_ _04345_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__mux2_1
XFILLER_44_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13708_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__xnor2_1
X_17476_ _09933_ _09936_ _10041_ vssd1 vssd1 vccd1 vccd1 _10042_ sky130_fd_sc_hd__a21oi_2
X_14688_ _07378_ _07413_ _06239_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__a21oi_1
XFILLER_204_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19215_ _02756_ vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__clkbuf_1
X_13639_ _06332_ _06331_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__xor2_1
X_16427_ _09069_ _09070_ _09071_ vssd1 vssd1 vccd1 vccd1 _09072_ sky130_fd_sc_hd__a21o_1
XFILLER_177_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16358_ _07967_ _08674_ _08034_ _08045_ vssd1 vssd1 vccd1 vccd1 _09003_ sky130_fd_sc_hd__or4_1
X_19146_ rbzero.spi_registers.new_other\[6\] _02712_ vssd1 vssd1 vccd1 vccd1 _02713_
+ sky130_fd_sc_hd__or2_1
XFILLER_173_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__04835_ _04835_ vssd1 vssd1 vccd1 vccd1 clknet_0__04835_ sky130_fd_sc_hd__clkbuf_16
XFILLER_146_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15309_ _07952_ _07953_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__and2_1
XFILLER_173_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16289_ _08908_ _08930_ _08931_ _08933_ vssd1 vssd1 vccd1 vccd1 _08934_ sky130_fd_sc_hd__and4_1
X_19077_ rbzero.pov.spi_buffer\[69\] rbzero.pov.ready_buffer\[69\] _02594_ vssd1 vssd1
+ vccd1 vccd1 _02671_ sky130_fd_sc_hd__mux2_1
XFILLER_161_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18028_ _01728_ _01729_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__xor2_1
XFILLER_172_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19979_ rbzero.pov.ready_buffer\[28\] _03252_ _03253_ rbzero.debug_overlay.facingY\[-3\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__o221a_1
XFILLER_80_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ clknet_leaf_49_i_clk _00592_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20754_ clknet_leaf_40_i_clk _00523_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[6\] sky130_fd_sc_hd__dfxtp_4
XFILLER_126_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20685_ clknet_leaf_65_i_clk _00469_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21306_ net227 _01075_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21237_ clknet_leaf_79_i_clk _01006_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21168_ clknet_leaf_92_i_clk _00937_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_172_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13990_ _06134_ _06677_ _06697_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__o21bai_1
X_21099_ net189 _00868_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ _05605_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__clkinv_2
XFILLER_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _08188_ _08239_ _08302_ _08304_ vssd1 vssd1 vccd1 vccd1 _08305_ sky130_fd_sc_hd__o31a_1
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _05561_ _05459_ _05608_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__o21a_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14611_ _07106_ _07337_ _07347_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__nand3_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _04598_ _04599_ _04218_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__mux2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _07970_ _08233_ _08234_ _08235_ vssd1 vssd1 vccd1 vccd1 _08236_ sky130_fd_sc_hd__o31ai_2
XFILLER_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ rbzero.wall_tracer.trackDistX\[-1\] rbzero.wall_tracer.stepDistX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _09898_ sky130_fd_sc_hd__nor2_1
XFILLER_199_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _07273_ _07278_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__or2b_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11754_ rbzero.tex_g0\[7\] rbzero.tex_g0\[6\] _04129_ vssd1 vssd1 vccd1 vccd1 _04532_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ rbzero.tex_g1\[5\] rbzero.tex_g1\[6\] _03691_ vssd1 vssd1 vccd1 vccd1 _03694_
+ sky130_fd_sc_hd__mux2_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ rbzero.wall_tracer.trackDistX\[-9\] _09836_ _05414_ vssd1 vssd1 vccd1 vccd1
+ _09837_ sky130_fd_sc_hd__mux2_1
X_14473_ _07204_ _07209_ _07154_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__a21oi_1
X_11685_ _04022_ _04440_ _04450_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__and3_2
X_16212_ _08227_ _08331_ _08856_ vssd1 vssd1 vccd1 vccd1 _08857_ sky130_fd_sc_hd__a21o_1
X_19000_ rbzero.pov.spi_buffer\[32\] rbzero.pov.ready_buffer\[32\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02631_ sky130_fd_sc_hd__mux2_1
X_13424_ _06119_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__clkbuf_4
XFILLER_186_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10636_ _03657_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__clkbuf_1
X_17192_ _09774_ _09776_ vssd1 vssd1 vccd1 vccd1 _09777_ sky130_fd_sc_hd__or2_1
X_16143_ _08266_ _08039_ _08040_ vssd1 vssd1 vccd1 vccd1 _08788_ sky130_fd_sc_hd__and3_1
X_13355_ _06036_ _06035_ _06030_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__a21bo_1
X_10567_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _03613_ vssd1 vssd1 vccd1 vccd1 _03621_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12306_ _04154_ _03477_ net20 vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__mux2_1
XFILLER_142_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16074_ _08692_ _08718_ vssd1 vssd1 vccd1 vccd1 _08719_ sky130_fd_sc_hd__xnor2_2
XFILLER_142_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13286_ _05973_ _06011_ _06009_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__o21a_1
X_10498_ rbzero.tex_r0\[40\] rbzero.tex_r0\[39\] _03580_ vssd1 vssd1 vccd1 vccd1 _03585_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15025_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__nand2_1
X_19902_ _07917_ _03141_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__nor2_1
X_12237_ net16 _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__or2_1
XFILLER_64_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19833_ rbzero.pov.ready_buffer\[62\] _07900_ _03146_ vssd1 vssd1 vccd1 vccd1 _03152_
+ sky130_fd_sc_hd__mux2_1
XFILLER_96_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12168_ _04021_ _04922_ _04905_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__and3_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11119_ _03910_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__clkbuf_1
X_19764_ _03110_ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12099_ _04862_ _04866_ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__o21a_1
X_16976_ _09614_ _09615_ vssd1 vssd1 vccd1 vccd1 _09616_ sky130_fd_sc_hd__nor2_1
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18715_ rbzero.wall_tracer.trackDistY\[-10\] rbzero.wall_tracer.stepDistY\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__nor2_1
Xinput6 i_gpout0_sel[4] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_8
X_15927_ _07945_ rbzero.wall_tracer.stepDistX\[-12\] _08135_ vssd1 vssd1 vccd1 vccd1
+ _08572_ sky130_fd_sc_hd__a21boi_4
X_19695_ _03074_ vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18646_ _02340_ _02341_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_0__03295_ _03295_ vssd1 vssd1 vccd1 vccd1 clknet_0__03295_ sky130_fd_sc_hd__clkbuf_16
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15858_ _08496_ _08502_ vssd1 vssd1 vccd1 vccd1 _08503_ sky130_fd_sc_hd__xor2_1
XFILLER_25_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14809_ _05884_ _07507_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__nor2_1
X_18577_ _09141_ _01475_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__nor2_1
X_15789_ _08432_ _08433_ vssd1 vssd1 vccd1 vccd1 _08434_ sky130_fd_sc_hd__xnor2_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17528_ _08202_ vssd1 vssd1 vccd1 vccd1 _10094_ sky130_fd_sc_hd__clkbuf_4
XFILLER_36_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17459_ _10023_ _10025_ vssd1 vssd1 vccd1 vccd1 _10026_ sky130_fd_sc_hd__xor2_4
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20095__129 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__inv_2
XFILLER_192_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20470_ rbzero.traced_texa\[-2\] rbzero.texV\[-2\] vssd1 vssd1 vccd1 vccd1 _03372_
+ sky130_fd_sc_hd__nor2_1
XFILLER_119_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19129_ _02699_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21022_ clknet_leaf_9_i_clk _00791_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_opt_2_0_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_2_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20806_ clknet_leaf_30_i_clk _00575_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20737_ clknet_leaf_81_i_clk _00506_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_196_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ _04211_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__buf_4
XFILLER_13_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20668_ clknet_leaf_61_i_clk _00452_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10421_ _03542_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20599_ _03462_ _03463_ rbzero.wall_tracer.rayAddendY\[-6\] _09762_ vssd1 vssd1 vccd1
+ vccd1 _01431_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13140_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__buf_2
XFILLER_109_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10352_ _03506_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _05804_ _05805_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__mux2_1
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ _04379_ _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__or2_1
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16830_ _09381_ _09348_ vssd1 vssd1 vccd1 vccd1 _09471_ sky130_fd_sc_hd__or2b_1
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16761_ _09393_ _09402_ vssd1 vssd1 vccd1 vccd1 _09403_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13973_ _06705_ _06709_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__nand2_1
XFILLER_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18500_ _02166_ _02197_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15712_ _08329_ _08356_ _08354_ vssd1 vssd1 vccd1 vccd1 _08357_ sky130_fd_sc_hd__o21ai_1
X_12924_ _05567_ _05660_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__nor2_1
XFILLER_111_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19480_ rbzero.wall_tracer.rayAddendY\[5\] _07855_ _02955_ _02960_ vssd1 vssd1 vccd1
+ vccd1 _00815_ sky130_fd_sc_hd__a211o_1
XFILLER_62_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16692_ _09331_ _09333_ vssd1 vssd1 vccd1 vccd1 _09335_ sky130_fd_sc_hd__nand2_1
XFILLER_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18431_ _02127_ _02129_ _09807_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a21oi_2
XFILLER_62_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15643_ _08285_ _08286_ _08287_ vssd1 vssd1 vccd1 vccd1 _08288_ sky130_fd_sc_hd__a21bo_1
X_12855_ rbzero.wall_tracer.visualWallDist\[-11\] rbzero.wall_tracer.rayAddendY\[-3\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__mux2_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _04217_ _04583_ _04123_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__o21a_1
X_18362_ _01960_ _01962_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__nor2_1
X_15574_ _08218_ _08208_ vssd1 vssd1 vccd1 vccd1 _08219_ sky130_fd_sc_hd__nand2_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ rbzero.wall_tracer.mapX\[5\] _05529_ _05414_ vssd1 vssd1 vccd1 vccd1 _05530_
+ sky130_fd_sc_hd__mux2_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14525_ _07077_ _07078_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__and2_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _09880_ _09881_ _09882_ vssd1 vssd1 vccd1 vccd1 _09883_ sky130_fd_sc_hd__and3_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ rbzero.debug_overlay.playerX\[-3\] _04463_ _04511_ _04513_ _04515_ vssd1
+ vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__a2111o_1
X_18293_ _01745_ _01988_ _01868_ _01869_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__a22oi_2
XFILLER_187_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14456_ _07191_ _07192_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__nor2_1
X_17244_ rbzero.wall_tracer.trackDistX\[-10\] rbzero.wall_tracer.stepDistX\[-10\]
+ vssd1 vssd1 vccd1 vccd1 _09821_ sky130_fd_sc_hd__or2_1
X_11668_ _03476_ _04441_ _04446_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a21bo_4
XFILLER_122_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13407_ _06131_ _06142_ _06143_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__a21o_1
X_10619_ rbzero.tex_g1\[46\] rbzero.tex_g1\[47\] _03647_ vssd1 vssd1 vccd1 vccd1 _03649_
+ sky130_fd_sc_hd__mux2_1
X_17175_ rbzero.traced_texa\[3\] _09770_ _09769_ net514 vssd1 vssd1 vccd1 vccd1 _00560_
+ sky130_fd_sc_hd__a22o_1
X_14387_ _07121_ _07123_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__xnor2_1
X_11599_ rbzero.tex_r1\[57\] _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__and3_1
XFILLER_183_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16126_ _07981_ _08042_ _08720_ vssd1 vssd1 vccd1 vccd1 _08771_ sky130_fd_sc_hd__or3_1
XFILLER_128_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13338_ _06069_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__nand2_1
XFILLER_116_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16057_ rbzero.wall_tracer.visualWallDist\[-11\] _04014_ _07990_ _07936_ vssd1 vssd1
+ vccd1 vccd1 _08702_ sky130_fd_sc_hd__and4_1
XFILLER_115_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13269_ _06004_ _06005_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__nand2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15008_ _07674_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_142_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19816_ net38 _03137_ _02708_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__o21ai_2
XFILLER_111_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03316_ clknet_0__03316_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03316_
+ sky130_fd_sc_hd__clkbuf_16
X_19747_ _03101_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16959_ _09597_ _09598_ vssd1 vssd1 vccd1 vccd1 _09600_ sky130_fd_sc_hd__and2_1
XFILLER_84_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19678_ _03065_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18629_ _02296_ _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__xnor2_1
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_197_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21640_ clknet_leaf_29_i_clk _01409_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21571_ net492 _01340_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_11 _07988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_22 _09781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_33 net24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20522_ rbzero.traced_texa\[6\] rbzero.texV\[6\] vssd1 vssd1 vccd1 vccd1 _03416_
+ sky130_fd_sc_hd__nor2_1
XANTENNA_44 _07549_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_55 net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_66 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_77 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20453_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 _03358_
+ sky130_fd_sc_hd__nand2_1
XFILLER_118_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21005_ clknet_leaf_11_i_clk _00774_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_153_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10970_ rbzero.tex_b1\[7\] rbzero.tex_b1\[8\] _03828_ vssd1 vssd1 vccd1 vccd1 _03833_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12640_ _05382_ _05384_ _05381_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__o21bai_1
XFILLER_102_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12571_ rbzero.wall_tracer.rayAddendY\[10\] rbzero.wall_tracer.rayAddendY\[9\] rbzero.debug_overlay.facingY\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__o21ai_1
XFILLER_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14310_ _07045_ _07046_ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__xor2_1
XFILLER_184_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11522_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _04213_ vssd1 vssd1 vccd1 vccd1 _04302_
+ sky130_fd_sc_hd__mux2_1
XFILLER_141_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15290_ _07933_ _07934_ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__nand2_1
XFILLER_200_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14241_ _06974_ _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__or2_1
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11453_ _04210_ _04220_ _04231_ _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__a211o_1
XFILLER_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10404_ _03533_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14172_ _06907_ _06908_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__nand2_1
X_11384_ rbzero.row_render.size\[1\] vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__inv_2
XFILLER_192_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13123_ _05648_ _05775_ _05788_ _05789_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__or4_1
XFILLER_152_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10335_ _03497_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18980_ _02620_ vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17931_ _10110_ _09693_ _01519_ _01633_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__o31ai_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__clkbuf_4
XFILLER_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ rbzero.tex_b1\[61\] rbzero.tex_b1\[60\] _04337_ vssd1 vssd1 vccd1 vccd1 _04780_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17862_ _01564_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__inv_2
XFILLER_79_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16813_ _09451_ _09453_ vssd1 vssd1 vccd1 vccd1 _09455_ sky130_fd_sc_hd__and2_1
X_17793_ _08188_ _09276_ _08493_ _08044_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__or4_1
XFILLER_94_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19532_ rbzero.debug_overlay.vplaneY\[-1\] _02987_ vssd1 vssd1 vccd1 vccd1 _03008_
+ sky130_fd_sc_hd__nor2_1
XFILLER_207_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16744_ _09268_ _09384_ _09385_ vssd1 vssd1 vccd1 vccd1 _09386_ sky130_fd_sc_hd__a21o_1
XFILLER_47_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13956_ _06679_ _06692_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__nor2_1
XFILLER_35_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19463_ _02942_ _02943_ _07676_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__o21ai_1
X_12907_ _05562_ _05566_ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__and3_1
XFILLER_207_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16675_ _09239_ _09317_ vssd1 vssd1 vccd1 vccd1 _09318_ sky130_fd_sc_hd__xnor2_1
X_13887_ _06201_ _06052_ _06623_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__and3_1
XFILLER_59_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20126__158 clknet_1_1__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__inv_2
XFILLER_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18414_ _02106_ _02107_ _02111_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__nand3_1
XFILLER_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _05569_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__and2_1
X_15626_ _07487_ _07455_ _07548_ _07551_ vssd1 vssd1 vccd1 vccd1 _08271_ sky130_fd_sc_hd__a22o_1
X_19394_ rbzero.debug_overlay.vplaneY\[0\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__nand2_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18345_ _02042_ _02043_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__and2_1
XFILLER_187_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _05506_ _05507_ _05504_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__a21o_1
X_15557_ _08199_ _08201_ vssd1 vssd1 vccd1 vccd1 _08202_ sky130_fd_sc_hd__nand2_4
XFILLER_30_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14508_ _07236_ _07243_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__nor2_1
X_18276_ _01973_ _01974_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__and2_1
X_15488_ _07460_ _08132_ _07933_ vssd1 vssd1 vccd1 vccd1 _08133_ sky130_fd_sc_hd__mux2_1
XFILLER_187_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput20 i_gpout3_sel[0] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_6
X_17227_ _09804_ _09805_ vssd1 vssd1 vccd1 vccd1 _09806_ sky130_fd_sc_hd__nor2_1
Xinput31 i_gpout4_sel[5] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__buf_4
X_14439_ _06689_ _06740_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__nor2_1
Xinput42 i_reg_mosi vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_16
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17158_ rbzero.traced_texa\[-11\] _09766_ _09767_ rbzero.wall_tracer.visualWallDist\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__a22o_1
XFILLER_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16109_ _08742_ _08752_ vssd1 vssd1 vccd1 vccd1 _08754_ sky130_fd_sc_hd__nor2_1
XFILLER_6_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17089_ _09726_ _09728_ vssd1 vssd1 vccd1 vccd1 _09729_ sky130_fd_sc_hd__xor2_2
XFILLER_171_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21623_ clknet_leaf_27_i_clk _01392_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21554_ net475 _01323_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20505_ rbzero.traced_texa\[3\] rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 _03402_
+ sky130_fd_sc_hd__nand2_1
XFILLER_166_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21485_ net406 _01254_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20436_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 _03344_
+ sky130_fd_sc_hd__and2_1
XFILLER_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19579__36 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__inv_2
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13810_ _06499_ _06465_ _06546_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__or3_1
X_14790_ _07459_ _07519_ _07521_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__and3_1
XFILLER_180_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13741_ _05946_ _05899_ _06007_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__or3_1
XFILLER_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10953_ rbzero.tex_b1\[15\] rbzero.tex_b1\[16\] _03817_ vssd1 vssd1 vccd1 vccd1 _03824_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16460_ _08360_ _09009_ vssd1 vssd1 vccd1 vccd1 _09104_ sky130_fd_sc_hd__nand2_1
X_13672_ _06041_ _06406_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__or2_1
XFILLER_189_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884_ rbzero.tex_b1\[48\] rbzero.tex_b1\[49\] _03784_ vssd1 vssd1 vccd1 vccd1 _03788_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15411_ _08043_ _08055_ vssd1 vssd1 vccd1 vccd1 _08056_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12623_ _05375_ _05376_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__nor2_1
XFILLER_188_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16391_ _09034_ _09035_ vssd1 vssd1 vccd1 vccd1 _09036_ sky130_fd_sc_hd__xor2_1
XFILLER_19_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18130_ _01829_ _01830_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15342_ rbzero.debug_overlay.playerX\[-8\] _05496_ _07986_ _05196_ vssd1 vssd1 vccd1
+ vccd1 _07987_ sky130_fd_sc_hd__a211o_1
XFILLER_40_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12554_ _05289_ _05295_ _05300_ _05307_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__and4_1
XFILLER_169_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11505_ rbzero.tex_r0\[3\] _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__and3_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18061_ _01760_ _01761_ _01756_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a21o_1
X_15273_ _07917_ rbzero.debug_overlay.playerY\[-5\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _07918_ sky130_fd_sc_hd__mux2_2
XFILLER_185_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12485_ rbzero.wall_tracer.trackDistX\[-9\] vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__03319_ clknet_0__03319_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03319_
+ sky130_fd_sc_hd__clkbuf_16
X_17012_ _09650_ _09651_ vssd1 vssd1 vccd1 vccd1 _09652_ sky130_fd_sc_hd__nor2_1
X_14224_ _06953_ _06960_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__xnor2_1
X_11436_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _04214_ vssd1 vssd1 vccd1 vccd1 _04216_
+ sky130_fd_sc_hd__mux2_1
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14155_ _06890_ _06891_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11367_ rbzero.row_render.size\[2\] vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__inv_2
XFILLER_152_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13106_ _05841_ _05842_ _05807_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__mux2_1
X_10318_ _03488_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_180_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14086_ _06802_ _06811_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__xnor2_1
X_18963_ _02611_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__clkbuf_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11298_ rbzero.traced_texVinit\[3\] rbzero.spi_registers.vshift\[0\] vssd1 vssd1
+ vccd1 vccd1 _04078_ sky130_fd_sc_hd__or2_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _08257_ _08044_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__nor2_1
XFILLER_152_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _05716_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__nor2_1
XFILLER_152_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18894_ _02560_ _02563_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__nor2_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17845_ _01441_ _01547_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__and2_1
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17776_ _07974_ _08427_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__nor2_1
X_14988_ _00008_ _07555_ _07664_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19515_ _02906_ rbzero.debug_overlay.vplaneY\[0\] vssd1 vssd1 vccd1 vccd1 _02993_
+ sky130_fd_sc_hd__and2_1
XFILLER_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16727_ _09368_ _08427_ vssd1 vssd1 vccd1 vccd1 _09369_ sky130_fd_sc_hd__nor2_1
XFILLER_93_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13939_ _06605_ _06611_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__and2_1
XFILLER_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19446_ _02927_ _02928_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__nand2_1
X_16658_ _09143_ _09140_ vssd1 vssd1 vccd1 vccd1 _09301_ sky130_fd_sc_hd__or2b_1
XFILLER_23_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_83_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15609_ _05193_ _08172_ _08174_ vssd1 vssd1 vccd1 vccd1 _08254_ sky130_fd_sc_hd__a21o_1
X_19377_ rbzero.debug_overlay.vplaneY\[-6\] _02849_ vssd1 vssd1 vccd1 vccd1 _02865_
+ sky130_fd_sc_hd__or2_1
XFILLER_176_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16589_ _09003_ _09006_ _09173_ vssd1 vssd1 vccd1 vccd1 _09232_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18328_ _10110_ _02026_ _01967_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__o21a_1
XFILLER_31_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18259_ _01953_ _01958_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_98_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_163_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21270_ clknet_leaf_93_i_clk _01039_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-7\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_156_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_21_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_143_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__buf_1
XFILLER_100_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_36_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20109__142 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__inv_2
X_20985_ clknet_leaf_11_i_clk _00754_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20261__279 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__inv_2
XFILLER_81_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21606_ net147 _01375_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21537_ net458 _01306_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12270_ _04891_ _04992_ _04890_ _04892_ _05024_ _05021_ vssd1 vssd1 vccd1 vccd1 _05039_
+ sky130_fd_sc_hd__mux4_1
XFILLER_175_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21468_ net389 _01237_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ gpout0.hpos\[5\] gpout0.hpos\[4\] gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1
+ _04008_ sky130_fd_sc_hd__and3_1
X_20419_ _03325_ _03328_ _03329_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__nand3b_1
XFILLER_150_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20155__184 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__inv_2
X_21399_ net320 _01168_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11152_ rbzero.debug_overlay.playerX\[5\] rbzero.wall_tracer.mapX\[5\] vssd1 vssd1
+ vccd1 vccd1 _03941_ sky130_fd_sc_hd__nand2_1
XFILLER_108_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11083_ rbzero.tex_b0\[18\] rbzero.tex_b0\[17\] _03887_ vssd1 vssd1 vccd1 vccd1 _03892_
+ sky130_fd_sc_hd__mux2_1
X_15960_ _08587_ _08604_ vssd1 vssd1 vccd1 vccd1 _08605_ sky130_fd_sc_hd__xor2_2
XFILLER_1_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14911_ _07591_ _07614_ _07615_ _04039_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__o211a_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _08505_ _08489_ vssd1 vssd1 vccd1 vccd1 _08536_ sky130_fd_sc_hd__xnor2_1
XFILLER_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17630_ _10042_ _10194_ vssd1 vssd1 vccd1 vccd1 _10195_ sky130_fd_sc_hd__xor2_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14842_ _07459_ _07453_ _07468_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__o21bai_4
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17561_ _10125_ _10126_ vssd1 vssd1 vccd1 vccd1 _10127_ sky130_fd_sc_hd__or2_1
XFILLER_91_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11985_ rbzero.tex_b1\[11\] _04221_ _04222_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__and3_1
XFILLER_17_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14773_ _07477_ _07476_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__nor2_1
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19300_ rbzero.spi_registers.new_other\[4\] rbzero.spi_registers.spi_buffer\[4\]
+ _02801_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__mux2_1
X_16512_ _09153_ _09155_ vssd1 vssd1 vccd1 vccd1 _09156_ sky130_fd_sc_hd__xor2_2
XFILLER_16_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13724_ _06391_ _06419_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10936_ rbzero.tex_b1\[23\] rbzero.tex_b1\[24\] _03806_ vssd1 vssd1 vccd1 vccd1 _03815_
+ sky130_fd_sc_hd__mux2_1
X_17492_ _09245_ _09029_ _09165_ _09243_ vssd1 vssd1 vccd1 vccd1 _10058_ sky130_fd_sc_hd__o22ai_1
XFILLER_204_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20320__332 clknet_1_0__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__inv_2
XFILLER_17_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19231_ rbzero.spi_registers.new_vshift\[2\] _02763_ vssd1 vssd1 vccd1 vccd1 _02767_
+ sky130_fd_sc_hd__or2_1
XFILLER_108_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16443_ _09059_ _08547_ vssd1 vssd1 vccd1 vccd1 _09087_ sky130_fd_sc_hd__and2b_1
XFILLER_32_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10867_ rbzero.tex_b1\[56\] rbzero.tex_b1\[57\] _03773_ vssd1 vssd1 vccd1 vccd1 _03779_
+ sky130_fd_sc_hd__mux2_1
X_13655_ _06351_ _06369_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__xor2_1
XFILLER_20_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19162_ rbzero.othery\[1\] _02710_ _02720_ _02722_ vssd1 vssd1 vccd1 vccd1 _00735_
+ sky130_fd_sc_hd__o211a_1
X_12606_ _05358_ _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__xnor2_2
X_16374_ _09008_ _09018_ vssd1 vssd1 vccd1 vccd1 _09019_ sky130_fd_sc_hd__xor2_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _06305_ _06321_ _06322_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ rbzero.tex_g0\[26\] rbzero.tex_g0\[25\] _03740_ vssd1 vssd1 vccd1 vccd1 _03743_
+ sky130_fd_sc_hd__mux2_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18113_ _01805_ _01806_ _01813_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a21oi_1
X_12537_ rbzero.debug_overlay.facingY\[-8\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__xor2_2
X_15325_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__buf_6
XFILLER_129_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19093_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.spi_buffer\[1\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__mux2_1
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ _01744_ _01745_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__xnor2_1
XFILLER_145_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12468_ _05220_ rbzero.wall_tracer.trackDistX\[6\] rbzero.wall_tracer.trackDistY\[5\]
+ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a2bb2o_1
X_15256_ rbzero.debug_overlay.playerX\[-6\] vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__inv_2
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11419_ gpout0.hpos\[6\] _04184_ _04182_ gpout0.hpos\[7\] _04198_ vssd1 vssd1 vccd1
+ vccd1 _04199_ sky130_fd_sc_hd__o221a_1
X_14207_ _06942_ _06943_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__nand2_1
X_15187_ _07829_ _07832_ _07840_ vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__o21bai_1
X_12399_ _04006_ _03475_ _04992_ _04892_ _05143_ net34 vssd1 vssd1 vccd1 vccd1 _05166_
+ sky130_fd_sc_hd__mux4_1
XFILLER_126_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14138_ _06860_ _06874_ _06872_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__a21o_1
XFILLER_152_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19995_ rbzero.pov.ready_buffer\[21\] _03252_ _03253_ _07821_ _03254_ vssd1 vssd1
+ vccd1 vccd1 _01036_ sky130_fd_sc_hd__o221a_1
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18946_ _02602_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__clkbuf_1
X_14069_ _06805_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__and3b_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18877_ _02549_ _02316_ rbzero.wall_tracer.trackDistY\[10\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00623_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17828_ _01530_ _01531_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__nor2_1
XFILLER_95_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17759_ _01462_ _09029_ _09165_ _09526_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__o22a_1
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20770_ clknet_leaf_43_i_clk _00539_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.texu\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19429_ _04471_ rbzero.debug_overlay.vplaneY\[-7\] _02910_ _02911_ vssd1 vssd1 vccd1
+ vccd1 _02913_ sky130_fd_sc_hd__or4_1
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21322_ net243 _01091_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21253_ clknet_leaf_85_i_clk _01022_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_190_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21184_ clknet_leaf_74_i_clk _00953_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11770_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _04341_ vssd1 vssd1 vccd1 vccd1 _04548_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20968_ clknet_leaf_7_i_clk _00737_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10721_ rbzero.tex_g0\[62\] rbzero.tex_g0\[61\] _03624_ vssd1 vssd1 vccd1 vccd1 _03702_
+ sky130_fd_sc_hd__mux2_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20899_ clknet_leaf_85_i_clk _00668_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ _06115_ _06176_ _06085_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__and3_1
X_10652_ rbzero.tex_g1\[30\] rbzero.tex_g1\[31\] _03658_ vssd1 vssd1 vccd1 vccd1 _03666_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13371_ _06097_ _06098_ _06106_ _06107_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__a31o_1
X_10583_ _03629_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12322_ net31 vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__inv_2
X_15110_ _07756_ _07761_ _07762_ _07768_ vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__a31o_1
X_16090_ _08570_ _08579_ _08571_ vssd1 vssd1 vccd1 vccd1 _08735_ sky130_fd_sc_hd__o21a_1
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15041_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__or2_1
X_12253_ _05021_ _04666_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__nand2_1
XFILLER_5_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11204_ _03988_ _03989_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__or3b_1
X_12184_ net13 _04953_ _04954_ _04922_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__a22o_1
XFILLER_69_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18800_ _02482_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__inv_2
X_11135_ rbzero.map_rom.f3 vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__clkinv_2
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19780_ rbzero.pov.spi_buffer\[63\] rbzero.pov.spi_buffer\[64\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03119_ sky130_fd_sc_hd__mux2_1
X_16992_ _08335_ _09217_ _09489_ _09490_ vssd1 vssd1 vccd1 vccd1 _09632_ sky130_fd_sc_hd__o31a_1
XFILLER_27_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.stepDistY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__and2_1
X_11066_ rbzero.tex_b0\[26\] rbzero.tex_b0\[25\] _03876_ vssd1 vssd1 vccd1 vccd1 _03883_
+ sky130_fd_sc_hd__mux2_1
X_15943_ _08526_ _08528_ vssd1 vssd1 vccd1 vccd1 _08588_ sky130_fd_sc_hd__xnor2_2
XFILLER_27_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18662_ _02255_ _02357_ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__xnor2_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15874_ _08518_ vssd1 vssd1 vccd1 vccd1 _08519_ sky130_fd_sc_hd__buf_4
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17613_ rbzero.wall_tracer.trackDistX\[1\] _09817_ _10173_ _10178_ vssd1 vssd1 vccd1
+ vccd1 _00590_ sky130_fd_sc_hd__o22a_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825_ _07473_ _07527_ _07499_ _07376_ _05834_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__a32o_2
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18593_ _02163_ _02199_ _02289_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a21oi_1
XFILLER_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _09114_ vssd1 vssd1 vccd1 vccd1 _10110_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _07351_ _07361_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__nor2_1
XFILLER_205_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11968_ rbzero.tex_b1\[23\] rbzero.tex_b1\[22\] _04290_ vssd1 vssd1 vccd1 vccd1 _04743_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13707_ _05846_ _06009_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__or2_1
X_17475_ _08416_ _09704_ _09924_ _09922_ vssd1 vssd1 vccd1 vccd1 _10041_ sky130_fd_sc_hd__o31a_1
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10919_ _03646_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__clkbuf_4
XFILLER_205_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11899_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _04290_ vssd1 vssd1 vccd1 vccd1 _04675_
+ sky130_fd_sc_hd__mux2_1
X_14687_ _07106_ _07419_ _07420_ _07423_ _05742_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__a311oi_2
XFILLER_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19214_ _09753_ _02755_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__and2_1
X_16426_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerX\[-8\] _07895_
+ vssd1 vssd1 vccd1 vccd1 _09071_ sky130_fd_sc_hd__mux2_1
X_13638_ _06347_ _06373_ _06374_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__a21boi_2
XFILLER_60_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19145_ rbzero.spi_registers.got_new_other _02711_ vssd1 vssd1 vccd1 vccd1 _02712_
+ sky130_fd_sc_hd__nand2_2
X_16357_ _08289_ _08294_ _09001_ vssd1 vssd1 vccd1 vccd1 _09002_ sky130_fd_sc_hd__a21bo_1
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13569_ _06097_ _06098_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__and2_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15308_ rbzero.debug_overlay.playerY\[-5\] _07906_ rbzero.debug_overlay.playerY\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__o21ai_1
X_19076_ _02670_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__clkbuf_1
X_16288_ _08901_ _08932_ vssd1 vssd1 vccd1 vccd1 _08933_ sky130_fd_sc_hd__nor2_1
XFILLER_146_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18027_ _01592_ _01601_ _01599_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a21oi_1
X_15239_ rbzero.wall_tracer.rayAddendX\[11\] _07887_ vssd1 vssd1 vccd1 vccd1 _07888_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_172_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19978_ _03242_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__buf_2
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18929_ rbzero.spi_registers.spi_counter\[6\] _02589_ _02592_ vssd1 vssd1 vccd1 vccd1
+ _00632_ sky130_fd_sc_hd__a21oi_1
XFILLER_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20822_ clknet_leaf_49_i_clk _00591_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20753_ clknet_leaf_40_i_clk _00522_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20684_ clknet_leaf_64_i_clk _00468_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_206_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21305_ net226 _01074_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21236_ clknet_leaf_79_i_clk _01005_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21167_ clknet_leaf_91_i_clk _00936_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21098_ net188 _00867_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_74_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20049_ _04891_ _03281_ _04890_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__a21oi_1
X_20267__285 clknet_1_1__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__inv_2
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12940_ _05675_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__xor2_2
XFILLER_105_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _04030_ _05367_ _05368_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__a31o_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14610_ _07343_ _07344_ _07346_ _07107_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__o211ai_2
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ rbzero.tex_g1\[53\] rbzero.tex_g1\[52\] _04212_ vssd1 vssd1 vccd1 vccd1 _04599_
+ sky130_fd_sc_hd__mux2_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _07970_ _08222_ _08223_ _08002_ vssd1 vssd1 vccd1 vccd1 _08235_ sky130_fd_sc_hd__a31oi_4
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14541_ _07276_ _07277_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__nor2_1
XFILLER_92_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _04129_ vssd1 vssd1 vccd1 vccd1 _04531_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10704_ _03693_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__clkbuf_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17260_ _09812_ _09833_ _09834_ _09835_ vssd1 vssd1 vccd1 vccd1 _09836_ sky130_fd_sc_hd__o31ai_1
XFILLER_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14472_ _07148_ _07208_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__xnor2_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _04004_ _04438_ _04450_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__and3_2
XFILLER_144_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16211_ _08377_ _08054_ vssd1 vssd1 vccd1 vccd1 _08856_ sky130_fd_sc_hd__nor2_1
X_10635_ rbzero.tex_g1\[38\] rbzero.tex_g1\[39\] _03647_ vssd1 vssd1 vccd1 vccd1 _03657_
+ sky130_fd_sc_hd__mux2_1
X_13423_ _05983_ _06159_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__nor2_1
X_17191_ rbzero.wall_tracer.mapX\[5\] _05512_ _09775_ vssd1 vssd1 vccd1 vccd1 _09776_
+ sky130_fd_sc_hd__o21a_1
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16142_ _08782_ _08783_ _08786_ vssd1 vssd1 vccd1 vccd1 _08787_ sky130_fd_sc_hd__o21ai_2
X_13354_ _06051_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__xnor2_1
X_10566_ _03620_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12305_ net22 _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__or2_1
XFILLER_182_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13285_ _06014_ _06018_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__xor2_2
X_16073_ _08693_ _08717_ vssd1 vssd1 vccd1 vccd1 _08718_ sky130_fd_sc_hd__xor2_2
X_10497_ _03584_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _04813_ _04811_ _04006_ _03475_ _04961_ _04960_ vssd1 vssd1 vccd1 vccd1 _05006_
+ sky130_fd_sc_hd__mux4_1
X_15024_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] _07688_
+ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__a21oi_1
X_19901_ rbzero.debug_overlay.playerY\[-6\] _03198_ _03204_ _03157_ vssd1 vssd1 vccd1
+ vccd1 _00992_ sky130_fd_sc_hd__o211a_1
XFILLER_29_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19832_ _03139_ _03150_ _03151_ _02765_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__o211a_1
X_12167_ net41 net43 net8 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__mux2_1
XFILLER_116_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11118_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _03557_ vssd1 vssd1 vccd1 vccd1 _03910_
+ sky130_fd_sc_hd__mux2_1
X_19763_ rbzero.pov.spi_buffer\[55\] rbzero.pov.spi_buffer\[56\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03110_ sky130_fd_sc_hd__mux2_1
X_12098_ _04868_ _04851_ _04855_ _04869_ net7 vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a32o_1
X_16975_ _09514_ _09607_ _09613_ vssd1 vssd1 vccd1 vccd1 _09615_ sky130_fd_sc_hd__and3_1
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18714_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ _02403_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a21oi_1
X_15926_ _08109_ _08491_ vssd1 vssd1 vccd1 vccd1 _08571_ sky130_fd_sc_hd__or2_1
X_11049_ rbzero.tex_b0\[34\] rbzero.tex_b0\[33\] _03865_ vssd1 vssd1 vccd1 vccd1 _03874_
+ sky130_fd_sc_hd__mux2_1
X_19694_ rbzero.pov.spi_buffer\[22\] rbzero.pov.spi_buffer\[23\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03074_ sky130_fd_sc_hd__mux2_1
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 i_gpout0_sel[5] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_8
XFILLER_77_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18645_ _10094_ _09611_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__03294_ _03294_ vssd1 vssd1 vccd1 vccd1 clknet_0__03294_ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _08497_ _08501_ _08499_ vssd1 vssd1 vccd1 vccd1 _08502_ sky130_fd_sc_hd__a21boi_1
XFILLER_65_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14808_ _00004_ _07536_ _07537_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a21oi_1
XFILLER_92_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18576_ _08151_ _09138_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__nor2_1
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _08161_ _08165_ vssd1 vssd1 vccd1 vccd1 _08433_ sky130_fd_sc_hd__or2_1
XFILLER_33_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17527_ _08178_ _08202_ _08493_ _08044_ vssd1 vssd1 vccd1 vccd1 _10093_ sky130_fd_sc_hd__or4_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14739_ _07378_ _07360_ vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__and2_1
XFILLER_71_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17458_ _09474_ _09733_ _10024_ vssd1 vssd1 vccd1 vccd1 _10025_ sky130_fd_sc_hd__a21oi_4
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16409_ _08437_ vssd1 vssd1 vccd1 vccd1 _09054_ sky130_fd_sc_hd__inv_2
XFILLER_193_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17389_ _09673_ _09676_ vssd1 vssd1 vccd1 vccd1 _09956_ sky130_fd_sc_hd__nor2_1
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19128_ rbzero.spi_registers.ss_buffer\[1\] rbzero.spi_registers.ss_buffer\[0\] _05189_
+ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__mux2_1
XFILLER_199_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19059_ rbzero.pov.spi_buffer\[60\] rbzero.pov.ready_buffer\[60\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02662_ sky130_fd_sc_hd__mux2_1
XFILLER_105_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21021_ clknet_leaf_8_i_clk _00790_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20805_ clknet_leaf_31_i_clk _00574_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20736_ clknet_leaf_82_i_clk _00505_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_156_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20667_ clknet_leaf_62_i_clk _00451_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10420_ rbzero.tex_r1\[10\] rbzero.tex_r1\[11\] _03538_ vssd1 vssd1 vccd1 vccd1 _03542_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20598_ _02827_ _02836_ _02835_ _07830_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__a31o_1
XFILLER_104_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10351_ rbzero.tex_r1\[43\] rbzero.tex_r1\[44\] _03505_ vssd1 vssd1 vccd1 vccd1 _03506_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13070_ _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12021_ rbzero.tex_b1\[33\] rbzero.tex_b1\[32\] _04250_ vssd1 vssd1 vccd1 vccd1 _04796_
+ sky130_fd_sc_hd__mux2_1
XFILLER_105_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21219_ clknet_leaf_19_i_clk _00988_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16760_ _09400_ _09401_ vssd1 vssd1 vccd1 vccd1 _09402_ sky130_fd_sc_hd__nor2_1
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13972_ _05825_ _06708_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__nor2_1
XFILLER_111_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15711_ _08059_ vssd1 vssd1 vccd1 vccd1 _08356_ sky130_fd_sc_hd__buf_4
XFILLER_150_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12923_ _05659_ _05569_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__and2_1
XFILLER_207_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16691_ _09331_ _09333_ vssd1 vssd1 vccd1 vccd1 _09334_ sky130_fd_sc_hd__nor2_1
XFILLER_19_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18430_ _01799_ _02024_ _02025_ _02023_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a22o_1
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15642_ _07977_ _07913_ _07924_ _07995_ vssd1 vssd1 vccd1 vccd1 _08287_ sky130_fd_sc_hd__or4_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12854_ rbzero.wall_tracer.rayAddendX\[-4\] _05590_ _05560_ vssd1 vssd1 vccd1 vccd1
+ _05591_ sky130_fd_sc_hd__mux2_2
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18361_ _02058_ _02059_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__nor2_1
X_11805_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _04211_ vssd1 vssd1 vccd1 vccd1 _04583_
+ sky130_fd_sc_hd__mux2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _07566_ vssd1 vssd1 vccd1 vccd1 _08218_ sky130_fd_sc_hd__inv_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ rbzero.debug_overlay.playerX\[5\] _05528_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05529_ sky130_fd_sc_hd__mux2_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _09872_ _09875_ _09873_ vssd1 vssd1 vccd1 vccd1 _09882_ sky130_fd_sc_hd__o21ai_1
XFILLER_42_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14524_ _07237_ _07260_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__xnor2_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18292_ _01990_ _01991_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__xor2_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ rbzero.debug_overlay.playerX\[2\] _04451_ _04465_ rbzero.debug_overlay.playerX\[-1\]
+ _04514_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__a221o_1
XFILLER_109_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17243_ _05242_ _09781_ _09820_ vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__a21oi_1
X_14455_ _07187_ _07190_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__nor2_1
X_11667_ gpout0.hpos\[8\] _04442_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__nand2_1
XFILLER_128_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13406_ _06130_ _06129_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__and2b_1
X_10618_ _03648_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17174_ _07706_ vssd1 vssd1 vccd1 vccd1 _09770_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11598_ _04375_ _04376_ _04219_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__mux2_1
X_14386_ _06698_ _06760_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__nor2_1
XFILLER_128_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16125_ _08180_ _08042_ _08769_ vssd1 vssd1 vccd1 vccd1 _08770_ sky130_fd_sc_hd__o21a_1
XFILLER_128_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10549_ _03611_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13337_ _06070_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__xor2_2
XFILLER_183_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16056_ _08644_ _08645_ vssd1 vssd1 vccd1 vccd1 _08701_ sky130_fd_sc_hd__xnor2_2
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13268_ _05983_ _05982_ _06003_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15007_ rbzero.wall_tracer.stepDistX\[10\] _07586_ _05201_ vssd1 vssd1 vccd1 vccd1
+ _07674_ sky130_fd_sc_hd__mux2_1
XFILLER_29_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12219_ gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__buf_2
XFILLER_123_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13199_ _05931_ _05903_ _05935_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19815_ _03136_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__buf_2
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03315_ clknet_0__03315_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03315_
+ sky130_fd_sc_hd__clkbuf_16
X_16958_ _09597_ _09598_ vssd1 vssd1 vccd1 vccd1 _09599_ sky130_fd_sc_hd__nor2_1
X_19746_ rbzero.pov.spi_buffer\[47\] rbzero.pov.spi_buffer\[48\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03101_ sky130_fd_sc_hd__mux2_1
XFILLER_77_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15909_ _08475_ _08553_ vssd1 vssd1 vccd1 vccd1 _08554_ sky130_fd_sc_hd__xor2_1
X_19677_ rbzero.pov.spi_buffer\[14\] rbzero.pov.spi_buffer\[15\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03065_ sky130_fd_sc_hd__mux2_1
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16889_ _08178_ _08111_ vssd1 vssd1 vccd1 vccd1 _09530_ sky130_fd_sc_hd__nor2_1
XFILLER_92_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18628_ _02288_ _02290_ _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__o21a_1
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18559_ _10239_ _09350_ _09481_ _10094_ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__o22a_1
XFILLER_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21570_ net491 _01339_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[21\] sky130_fd_sc_hd__dfxtp_1
X_20103__137 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__inv_2
XFILLER_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_12 _07988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20521_ rbzero.texV\[5\] _03327_ _03332_ _03415_ vssd1 vssd1 vccd1 vccd1 _01401_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_23 _09807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 _07916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_56 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_67 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_78 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20452_ rbzero.traced_texa\[-5\] rbzero.texV\[-5\] vssd1 vssd1 vccd1 vccd1 _03357_
+ sky130_fd_sc_hd__or2_1
XFILLER_193_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21004_ clknet_leaf_10_i_clk _00773_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20184__209 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__inv_2
XFILLER_101_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20379__386 clknet_1_1__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__inv_2
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _05288_ _05319_ _05320_ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__o211ai_2
XFILLER_93_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11521_ _04299_ _04300_ _04266_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__mux2_1
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20719_ clknet_leaf_72_i_clk _00009_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_20078__114 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__inv_2
XFILLER_196_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11452_ _04119_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__buf_4
X_14240_ _06844_ _06973_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__nor2_1
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10403_ rbzero.tex_r1\[18\] rbzero.tex_r1\[19\] _03527_ vssd1 vssd1 vccd1 vccd1 _03533_
+ sky130_fd_sc_hd__mux2_1
X_14171_ _06887_ _06901_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__xor2_1
X_11383_ gpout0.hpos\[1\] vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__clkbuf_4
XFILLER_124_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10334_ rbzero.tex_r1\[51\] rbzero.tex_r1\[52\] _03494_ vssd1 vssd1 vccd1 vccd1 _03497_
+ sky130_fd_sc_hd__mux2_1
X_13122_ _05857_ _05858_ _05807_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__mux2_1
XFILLER_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17930_ _01514_ _01518_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__nand2_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _05775_ _05788_ _05789_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__or3_1
XFILLER_106_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12004_ rbzero.tex_b1\[63\] rbzero.tex_b1\[62\] _04337_ vssd1 vssd1 vccd1 vccd1 _04779_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17861_ _09249_ _10200_ _01458_ _01460_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__o22a_1
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16812_ _09451_ _09453_ vssd1 vssd1 vccd1 vccd1 _09454_ sky130_fd_sc_hd__nor2_1
XFILLER_113_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17792_ _10257_ _10263_ _01495_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__a21oi_2
XFILLER_120_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19531_ rbzero.wall_tracer.rayAddendY\[9\] _07718_ _07831_ _03005_ _03007_ vssd1
+ vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__o221a_1
X_16743_ _09269_ _09273_ vssd1 vssd1 vccd1 vccd1 _09385_ sky130_fd_sc_hd__and2_1
X_13955_ _06680_ _06672_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__nor2_1
XFILLER_4_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19462_ _02942_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__and2_1
X_12906_ _05610_ _05612_ _05615_ _05601_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__a211o_1
X_16674_ _09315_ _09316_ vssd1 vssd1 vccd1 vccd1 _09317_ sky130_fd_sc_hd__nor2_1
XFILLER_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _05974_ _05983_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__nand2_1
XFILLER_62_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18413_ _02106_ _02107_ _02111_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__a21o_1
XFILLER_146_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _07551_ vssd1 vssd1 vccd1 vccd1 _08270_ sky130_fd_sc_hd__inv_2
X_19393_ rbzero.debug_overlay.vplaneY\[0\] rbzero.wall_tracer.rayAddendY\[0\] vssd1
+ vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__or2_1
X_12837_ _05563_ _05573_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__nand2_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ _09141_ _01620_ _02041_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__o21ai_1
XFILLER_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15556_ _08002_ _08200_ _07945_ vssd1 vssd1 vccd1 vccd1 _08201_ sky130_fd_sc_hd__a21oi_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12768_ _05511_ _05513_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__or2b_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14507_ _07236_ _07243_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__nand2_1
X_18275_ _01973_ _01974_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__nor2_1
XFILLER_187_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11719_ rbzero.debug_overlay.playerY\[-5\] _04454_ _04458_ rbzero.debug_overlay.playerY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__a22o_1
X_15487_ rbzero.wall_tracer.rayAddendY\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] _07893_
+ vssd1 vssd1 vccd1 vccd1 _08132_ sky130_fd_sc_hd__mux2_1
X_12699_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[10\] vssd1
+ vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__xnor2_4
X_17226_ _08939_ _08850_ _08936_ vssd1 vssd1 vccd1 vccd1 _09805_ sky130_fd_sc_hd__and3_1
XFILLER_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput10 i_gpout1_sel[2] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_8
X_14438_ _07172_ _07174_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__xnor2_1
XFILLER_175_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput21 i_gpout3_sel[1] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_6
Xinput32 i_gpout5_sel[0] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_4
Xinput43 i_reg_sclk vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_8
X_17157_ rbzero.traced_texa\[-12\] _09766_ _09767_ rbzero.wall_tracer.visualWallDist\[-12\]
+ vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__a22o_1
X_14369_ _05931_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__buf_2
XFILLER_183_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16108_ _08742_ _08752_ vssd1 vssd1 vccd1 vccd1 _08753_ sky130_fd_sc_hd__xor2_1
XFILLER_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17088_ _09517_ _09582_ _09727_ vssd1 vssd1 vccd1 vccd1 _09728_ sky130_fd_sc_hd__a21oi_2
XFILLER_196_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16039_ _07958_ _08491_ vssd1 vssd1 vccd1 vccd1 _08684_ sky130_fd_sc_hd__or2_1
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19729_ _03047_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21622_ clknet_leaf_74_i_clk _01391_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21553_ net474 _01322_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20504_ rbzero.traced_texa\[3\] rbzero.texV\[3\] vssd1 vssd1 vccd1 vccd1 _03401_
+ sky130_fd_sc_hd__or2_1
XFILLER_194_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21484_ net405 _01253_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20435_ rbzero.traced_texa\[-8\] rbzero.texV\[-8\] vssd1 vssd1 vccd1 vccd1 _03343_
+ sky130_fd_sc_hd__nor2_1
XFILLER_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13740_ _05944_ _06016_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__nor2_1
X_10952_ _03823_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_189_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13671_ _06061_ _06407_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__nand2_1
X_10883_ _03787_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15410_ _08047_ _08054_ vssd1 vssd1 vccd1 vccd1 _08055_ sky130_fd_sc_hd__nor2_1
XFILLER_188_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ _03942_ _05374_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__nor2_1
X_16390_ _08062_ _08425_ vssd1 vssd1 vccd1 vccd1 _09035_ sky130_fd_sc_hd__nor2_1
XFILLER_19_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15341_ _05495_ _07985_ vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__nor2_1
XFILLER_19_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12553_ _05303_ _05306_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__and2_1
XFILLER_169_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18060_ _01756_ _01760_ _01761_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__nand3_1
X_11504_ _04282_ _04283_ _04226_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__mux2_1
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15272_ rbzero.debug_overlay.playerY\[-5\] _07906_ vssd1 vssd1 vccd1 vccd1 _07917_
+ sky130_fd_sc_hd__xor2_1
XFILLER_156_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03318_ clknet_0__03318_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03318_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12484_ rbzero.wall_tracer.trackDistX\[-8\] vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__inv_2
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17011_ _09647_ _09649_ vssd1 vssd1 vccd1 vccd1 _09651_ sky130_fd_sc_hd__and2_1
X_14223_ _06958_ _06959_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__and2b_1
X_11435_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _04214_ vssd1 vssd1 vccd1 vccd1 _04215_
+ sky130_fd_sc_hd__mux2_1
XFILLER_138_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11366_ _04137_ _04139_ _04140_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__or4_1
X_14154_ _06666_ _06672_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__nor2_1
XFILLER_99_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10317_ rbzero.tex_r1\[59\] rbzero.tex_r1\[60\] _03483_ vssd1 vssd1 vccd1 vccd1 _03488_
+ sky130_fd_sc_hd__mux2_1
X_13105_ _05690_ _05681_ _05791_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__mux2_1
XFILLER_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_2_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14085_ _06687_ _06694_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__xor2_1
X_18962_ rbzero.pov.spi_buffer\[14\] rbzero.pov.ready_buffer\[14\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02611_ sky130_fd_sc_hd__mux2_1
X_11297_ rbzero.texV\[4\] _04076_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__xor2_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20132__163 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__inv_2
X_17913_ _08242_ _09129_ _08129_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__a21oi_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _05598_ _05717_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__xnor2_2
XFILLER_156_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18893_ _02562_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__inv_2
XFILLER_152_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17844_ _01441_ _01547_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__nor2_1
XFILLER_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17775_ _01477_ _01478_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__nand2_1
X_14987_ rbzero.wall_tracer.stepDistX\[0\] _07650_ vssd1 vssd1 vccd1 vccd1 _07664_
+ sky130_fd_sc_hd__nor2_1
XFILLER_187_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16726_ _08823_ vssd1 vssd1 vccd1 vccd1 _09368_ sky130_fd_sc_hd__buf_2
X_19514_ _02990_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__nor2_1
X_13938_ _06240_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__clkbuf_4
XFILLER_170_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19445_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.debug_overlay.vplaneY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__nand2_1
XFILLER_179_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16657_ _09297_ _09298_ _09282_ vssd1 vssd1 vccd1 vccd1 _09300_ sky130_fd_sc_hd__a21o_1
XFILLER_23_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13869_ _06548_ _06549_ _06551_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__or3_1
Xclkbuf_0__03045_ _03045_ vssd1 vssd1 vccd1 vccd1 clknet_0__03045_ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15608_ _08183_ _08185_ _07598_ _08002_ _05208_ vssd1 vssd1 vccd1 vccd1 _08253_ sky130_fd_sc_hd__a2111o_1
X_19376_ _02862_ _02863_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16588_ _09223_ _09230_ vssd1 vssd1 vccd1 vccd1 _09231_ sky130_fd_sc_hd__xnor2_1
XFILLER_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18327_ _10134_ _01878_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__nand2_1
XFILLER_176_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _07894_ _05335_ vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__nor2_1
XFILLER_188_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18258_ _01956_ _01957_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__xor2_1
XFILLER_176_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ rbzero.wall_tracer.mapX\[8\] _05525_ _09790_ vssd1 vssd1 vccd1 vccd1 _09791_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_191_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18189_ _01887_ _01888_ _01889_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__nand3_1
XFILLER_191_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20215__238 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__inv_2
XFILLER_143_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ clknet_leaf_9_i_clk _00753_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19584__40 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__inv_2
XFILLER_129_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21605_ net146 _01374_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21536_ net457 _01305_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_103_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21467_ net388 _01236_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11220_ _04004_ _04005_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__o21ai_1
XFILLER_153_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20418_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 _03329_
+ sky130_fd_sc_hd__nand2_1
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21398_ net319 _01167_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ rbzero.debug_overlay.playerX\[5\] rbzero.wall_tracer.mapX\[5\] vssd1 vssd1
+ vccd1 vccd1 _03940_ sky130_fd_sc_hd__or2_1
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20349_ clknet_1_0__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__buf_1
XFILLER_134_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _03891_ vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14910_ rbzero.wall_tracer.visualWallDist\[-4\] _07595_ vssd1 vssd1 vccd1 vccd1 _07615_
+ sky130_fd_sc_hd__or2_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _08513_ _08534_ vssd1 vssd1 vccd1 vccd1 _08535_ sky130_fd_sc_hd__xor2_1
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ _07563_ vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__clkbuf_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _09700_ _09998_ vssd1 vssd1 vccd1 vccd1 _10126_ sky130_fd_sc_hd__and2_1
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14772_ _05814_ _07504_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__or2_1
X_11984_ rbzero.tex_b1\[9\] rbzero.tex_b1\[8\] _04263_ vssd1 vssd1 vccd1 vccd1 _04759_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16511_ _08998_ _09021_ _09154_ vssd1 vssd1 vccd1 vccd1 _09155_ sky130_fd_sc_hd__a21oi_2
XFILLER_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13723_ _06436_ _06459_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__or2b_1
XFILLER_204_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17491_ _10055_ _10056_ vssd1 vssd1 vccd1 vccd1 _10057_ sky130_fd_sc_hd__xnor2_1
XFILLER_17_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10935_ _03814_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20162__189 clknet_1_0__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__inv_2
X_19230_ rbzero.spi_registers.vshift\[1\] _02762_ _02766_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00759_ sky130_fd_sc_hd__o211a_1
XFILLER_140_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16442_ _09083_ _09084_ _09086_ _07642_ vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__o211a_1
XFILLER_140_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13654_ _06388_ _06390_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__and2_1
XFILLER_95_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10866_ _03778_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _05290_ _05293_ _05294_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__a21o_1
X_19161_ _02721_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__buf_2
X_16373_ _09016_ _09017_ vssd1 vssd1 vccd1 vccd1 _09018_ sky130_fd_sc_hd__nor2_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13585_ _06308_ _06320_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__and2b_1
XFILLER_157_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10797_ _03742_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__clkbuf_1
X_18112_ _01811_ _01812_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__nand2_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _07944_ _07968_ vssd1 vssd1 vccd1 vccd1 _07969_ sky130_fd_sc_hd__xor2_1
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19092_ _02679_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__clkbuf_1
X_12536_ rbzero.debug_overlay.facingY\[-7\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__or2_1
XFILLER_185_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18043_ _09292_ _09695_ _08802_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__a21oi_2
X_15255_ _07898_ _07899_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__nand2_1
X_12467_ rbzero.wall_tracer.trackDistX\[5\] vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__inv_2
XFILLER_32_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14206_ _06934_ _06939_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__xor2_1
XFILLER_67_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11418_ _04004_ _04186_ _04184_ gpout0.hpos\[6\] _04197_ vssd1 vssd1 vccd1 vccd1
+ _04198_ sky130_fd_sc_hd__a221o_1
XFILLER_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15186_ rbzero.wall_tracer.rayAddendX\[6\] _07695_ _07839_ _03913_ vssd1 vssd1 vccd1
+ vccd1 _07840_ sky130_fd_sc_hd__a22o_1
X_12398_ _05153_ _05149_ _05154_ _05164_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__o31a_1
XFILLER_141_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14137_ _06872_ _06873_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__and2b_1
X_11349_ _04128_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__buf_4
XFILLER_28_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19994_ rbzero.pov.ready_buffer\[20\] _03252_ _03253_ _07742_ _03254_ vssd1 vssd1
+ vccd1 vccd1 _01035_ sky130_fd_sc_hd__o221a_1
XFILLER_4_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18945_ rbzero.pov.spi_buffer\[6\] rbzero.pov.ready_buffer\[6\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02602_ sky130_fd_sc_hd__mux2_1
X_14068_ _06009_ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__buf_2
XFILLER_140_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13019_ _05736_ _05735_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__or2_1
XFILLER_79_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18876_ _05532_ _02548_ _02406_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__o21a_1
XFILLER_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17827_ _10264_ _10272_ _10271_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__a21oi_1
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17758_ _09522_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__buf_2
X_16709_ _05210_ _09350_ vssd1 vssd1 vccd1 vccd1 _09351_ sky130_fd_sc_hd__or2_1
X_17689_ _10235_ _10253_ vssd1 vssd1 vccd1 vccd1 _10254_ sky130_fd_sc_hd__xor2_2
XFILLER_63_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19428_ _04471_ rbzero.debug_overlay.vplaneY\[-7\] _02910_ _02911_ vssd1 vssd1 vccd1
+ vccd1 _02912_ sky130_fd_sc_hd__o22ai_1
XFILLER_50_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19359_ rbzero.wall_tracer.rayAddendY\[-4\] _00013_ _02845_ _02848_ vssd1 vssd1 vccd1
+ vccd1 _00806_ sky130_fd_sc_hd__o22a_1
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21321_ net242 _01090_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20139__169 clknet_1_0__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__inv_2
XFILLER_135_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21252_ clknet_leaf_87_i_clk _01021_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_191_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21183_ clknet_leaf_18_i_clk _00952_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19636__88 clknet_1_0__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__inv_2
XFILLER_131_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ clknet_leaf_8_i_clk _00736_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_867 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10720_ _03701_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ clknet_leaf_68_i_clk _00667_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_158_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10651_ _03665_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10582_ rbzero.tex_g1\[63\] net47 _03549_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__mux2_1
X_13370_ _06102_ _06105_ _06099_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__a21oi_1
XFILLER_186_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ _05087_ net61 _05088_ net30 vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__o211a_1
XFILLER_139_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21519_ net440 _01288_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15040_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__nand2_1
X_12252_ net20 vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__buf_2
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20350__359 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__inv_2
XFILLER_135_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11203_ rbzero.map_rom.f3 rbzero.map_rom.d6 _03990_ _03991_ vssd1 vssd1 vccd1 vccd1
+ _03992_ sky130_fd_sc_hd__o211a_1
X_12183_ net11 net10 _04904_ _04867_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__and4b_1
XFILLER_150_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11134_ rbzero.debug_overlay.playerX\[0\] _03919_ rbzero.map_rom.i_row\[4\] _03920_
+ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__a221o_1
X_16991_ _09627_ _09630_ vssd1 vssd1 vccd1 vccd1 _09631_ sky130_fd_sc_hd__xnor2_1
XFILLER_122_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_82_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18730_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.stepDistY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__nor2_1
X_11065_ _03882_ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__clkbuf_1
X_15942_ _08531_ _08532_ vssd1 vssd1 vccd1 vccd1 _08587_ sky130_fd_sc_hd__xnor2_2
XFILLER_88_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18661_ _02355_ _02356_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__nand2_1
XFILLER_95_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ _05195_ _08226_ vssd1 vssd1 vccd1 vccd1 _08518_ sky130_fd_sc_hd__or2_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824_ _00004_ _07549_ _07550_ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__a21oi_1
X_17612_ _09889_ _10176_ _10177_ _09780_ vssd1 vssd1 vccd1 vccd1 _10178_ sky130_fd_sc_hd__a31o_1
X_18592_ _02161_ _02162_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__nor2_1
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_97_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20244__264 clknet_1_0__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__inv_2
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17543_ _10090_ _10108_ vssd1 vssd1 vccd1 vccd1 _10109_ sky130_fd_sc_hd__xor2_2
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14755_ _07107_ _07349_ _07337_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__a21bo_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11967_ rbzero.tex_b1\[21\] rbzero.tex_b1\[20\] _04356_ vssd1 vssd1 vccd1 vccd1 _04742_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_205_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13706_ _05823_ _05909_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__or2_1
X_17474_ _09954_ _09919_ vssd1 vssd1 vccd1 vccd1 _10040_ sky130_fd_sc_hd__or2b_1
X_10918_ _03805_ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_20_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_14686_ _05779_ _07337_ _07347_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__and3_1
X_11898_ _04247_ _04671_ _04672_ _04673_ _04229_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__o221a_1
XFILLER_177_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19213_ rbzero.spi_registers.new_floor\[2\] rbzero.color_floor\[2\] _02751_ vssd1
+ vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__mux2_1
X_16425_ rbzero.debug_overlay.playerY\[-9\] rbzero.debug_overlay.playerX\[-9\] _07894_
+ vssd1 vssd1 vccd1 vccd1 _09070_ sky130_fd_sc_hd__mux2_1
XFILLER_204_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13637_ _06372_ _06349_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__or2b_1
X_10849_ _03769_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19144_ _02708_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__clkbuf_4
X_16356_ _08295_ _08288_ vssd1 vssd1 vccd1 vccd1 _09001_ sky130_fd_sc_hd__or2b_1
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13568_ _06291_ _06298_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__xor2_2
XFILLER_9_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15307_ rbzero.debug_overlay.playerY\[-4\] rbzero.debug_overlay.playerY\[-5\] _07906_
+ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__or3_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19075_ rbzero.pov.spi_buffer\[68\] rbzero.pov.ready_buffer\[68\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02670_ sky130_fd_sc_hd__mux2_1
X_12519_ _05261_ _05259_ _05256_ _05273_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__o211ai_1
XFILLER_200_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_35_i_clk clknet_opt_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_160_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16287_ _08900_ _08885_ _08888_ vssd1 vssd1 vccd1 vccd1 _08932_ sky130_fd_sc_hd__and3_1
XFILLER_145_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13499_ _05752_ _06153_ _06207_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__and3_1
XFILLER_69_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18026_ _01726_ _01727_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__nand2_1
X_15238_ _07885_ _07821_ _07886_ vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__mux2_1
XFILLER_145_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _07819_ _07822_ _07818_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__a21o_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19977_ _03239_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__clkbuf_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18928_ rbzero.spi_registers.spi_counter\[6\] _02589_ _02557_ vssd1 vssd1 vccd1 vccd1
+ _02592_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18859_ _02530_ _02531_ _02532_ _05203_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__o31a_1
XFILLER_131_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19641__91 clknet_1_0__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__inv_2
XFILLER_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20821_ clknet_leaf_48_i_clk _00590_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20752_ clknet_leaf_36_i_clk _00521_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20683_ clknet_leaf_65_i_clk _00467_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21304_ net225 _01073_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_152_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21235_ clknet_leaf_91_i_clk _01004_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21166_ clknet_leaf_89_i_clk _00935_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21097_ net187 _00866_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20048_ _04891_ _03281_ _03284_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__o21ba_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12870_ rbzero.wall_tracer.visualWallDist\[0\] _05571_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05607_ sky130_fd_sc_hd__a21o_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ rbzero.tex_g1\[55\] rbzero.tex_g1\[54\] _04212_ vssd1 vssd1 vccd1 vccd1 _04598_
+ sky130_fd_sc_hd__mux2_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _07274_ _07275_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__and2_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _04345_ _04527_ _04528_ _04529_ _04253_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__o221a_1
XFILLER_109_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10703_ rbzero.tex_g1\[6\] rbzero.tex_g1\[7\] _03691_ vssd1 vssd1 vccd1 vccd1 _03693_
+ sky130_fd_sc_hd__mux2_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14471_ _07206_ _07207_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__or2_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11683_ rbzero.debug_overlay.vplaneX\[-3\] vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__buf_4
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _08377_ _08329_ _08854_ vssd1 vssd1 vccd1 vccd1 _08855_ sky130_fd_sc_hd__or3b_1
X_13422_ _05995_ _06113_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__and2_1
XFILLER_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10634_ _03656_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__clkbuf_1
X_17190_ rbzero.wall_tracer.mapX\[5\] _05512_ _05527_ vssd1 vssd1 vccd1 vccd1 _09775_
+ sky130_fd_sc_hd__a21o_1
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16141_ _08594_ _08075_ _08784_ _08785_ vssd1 vssd1 vccd1 vccd1 _08786_ sky130_fd_sc_hd__o31a_1
XFILLER_139_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13353_ _06075_ _06089_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10565_ rbzero.tex_r0\[8\] rbzero.tex_r0\[7\] _03613_ vssd1 vssd1 vccd1 vccd1 _03620_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _04813_ _04811_ _04006_ _03475_ net20 net21 vssd1 vssd1 vccd1 vccd1 _05073_
+ sky130_fd_sc_hd__mux4_1
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16072_ _08695_ _08715_ _08716_ vssd1 vssd1 vccd1 vccd1 _08717_ sky130_fd_sc_hd__a21oi_2
X_13284_ _06001_ _06020_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__xnor2_1
X_10496_ rbzero.tex_r0\[41\] rbzero.tex_r0\[40\] _03580_ vssd1 vssd1 vccd1 vccd1 _03584_
+ sky130_fd_sc_hd__mux2_1
XFILLER_170_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15023_ _07685_ _07686_ _07687_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__and3b_1
X_19900_ rbzero.pov.ready_buffer\[47\] _02823_ _03193_ _03203_ vssd1 vssd1 vccd1 vccd1
+ _03204_ sky130_fd_sc_hd__a211o_1
X_12235_ _04154_ _03477_ _04966_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__mux2_1
XFILLER_107_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19831_ _08000_ _03143_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__nand2_1
X_12166_ net39 _04918_ _04936_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a21o_1
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11117_ _03909_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19762_ _03109_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__clkbuf_1
X_12097_ net6 vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__inv_2
X_16974_ _09514_ _09607_ _09613_ vssd1 vssd1 vccd1 vccd1 _09614_ sky130_fd_sc_hd__a21oi_4
X_18713_ _02405_ _09819_ rbzero.wall_tracer.trackDistY\[-11\] _02406_ vssd1 vssd1
+ vccd1 vccd1 _00602_ sky130_fd_sc_hd__o2bb2a_1
X_15925_ _08084_ vssd1 vssd1 vccd1 vccd1 _08570_ sky130_fd_sc_hd__buf_4
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11048_ _03873_ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__clkbuf_1
X_19693_ _03073_ vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__clkbuf_1
Xinput8 i_gpout1_sel[0] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_16
XFILLER_49_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20168__195 clknet_1_0__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__inv_2
XFILLER_65_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18644_ _02335_ _02339_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__xnor2_1
X_15856_ _08499_ _08500_ vssd1 vssd1 vccd1 vccd1 _08501_ sky130_fd_sc_hd__and2_1
Xclkbuf_0__03293_ _03293_ vssd1 vssd1 vccd1 vccd1 clknet_0__03293_ sky130_fd_sc_hd__clkbuf_16
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14807_ rbzero.wall_tracer.stepDistY\[-5\] _07461_ vssd1 vssd1 vccd1 vccd1 _07537_
+ sky130_fd_sc_hd__nor2_1
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18575_ _02146_ _02148_ _02145_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a21bo_1
X_15787_ _08430_ _08431_ vssd1 vssd1 vccd1 vccd1 _08432_ sky130_fd_sc_hd__nor2_1
XFILLER_75_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12999_ _05687_ _05719_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__or2_2
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17526_ _09975_ _09985_ _10091_ vssd1 vssd1 vccd1 vccd1 _10092_ sky130_fd_sc_hd__a21oi_2
X_14738_ _05844_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__buf_2
XFILLER_205_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17457_ _09730_ _09732_ vssd1 vssd1 vccd1 vccd1 _10024_ sky130_fd_sc_hd__nor2_1
XFILLER_33_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14669_ _07376_ _07392_ _07405_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__or3_1
XFILLER_60_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16408_ _09050_ _09052_ vssd1 vssd1 vccd1 vccd1 _09053_ sky130_fd_sc_hd__xor2_2
XFILLER_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17388_ _09919_ _09954_ vssd1 vssd1 vccd1 vccd1 _09955_ sky130_fd_sc_hd__xnor2_2
XFILLER_192_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16339_ _05194_ _08982_ _08983_ _08224_ vssd1 vssd1 vccd1 vccd1 _08984_ sky130_fd_sc_hd__a31o_1
X_19127_ _02698_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__clkbuf_1
XFILLER_158_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19058_ _02661_ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18009_ _01581_ _01585_ _01583_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__a21boi_1
XFILLER_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21020_ clknet_leaf_8_i_clk _00789_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20385__11 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__inv_2
XFILLER_167_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20804_ clknet_leaf_30_i_clk _00573_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20735_ clknet_leaf_82_i_clk _00504_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20666_ clknet_leaf_63_i_clk _00450_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_91_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20597_ _02827_ _02836_ _02835_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__a21oi_1
XFILLER_192_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _03482_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__clkbuf_4
XFILLER_137_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12020_ _04254_ _04790_ _04794_ _04371_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a211o_1
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21218_ clknet_leaf_19_i_clk _00987_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21149_ clknet_leaf_86_i_clk _00918_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13971_ _06707_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15710_ _08354_ _08329_ _08058_ vssd1 vssd1 vccd1 vccd1 _08355_ sky130_fd_sc_hd__or3_1
XFILLER_74_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12922_ _04001_ _05494_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__nand2_1
XFILLER_207_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16690_ _09332_ _07949_ _07895_ vssd1 vssd1 vccd1 vccd1 _09333_ sky130_fd_sc_hd__mux2_1
XFILLER_150_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15641_ _07959_ _07932_ vssd1 vssd1 vccd1 vccd1 _08286_ sky130_fd_sc_hd__nor2_1
XFILLER_46_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12853_ rbzero.wall_tracer.visualWallDist\[-12\] rbzero.wall_tracer.rayAddendY\[-4\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__mux2_1
XFILLER_74_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _02056_ _02057_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__and2_1
X_11804_ _04224_ _04581_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__or2_1
XFILLER_15_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _08002_ rbzero.wall_tracer.stepDistY\[4\] vssd1 vssd1 vccd1 vccd1 _08217_
+ sky130_fd_sc_hd__and2_1
X_12784_ _05526_ _05527_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__xnor2_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ rbzero.wall_tracer.trackDistX\[-3\] rbzero.wall_tracer.stepDistX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _09881_ sky130_fd_sc_hd__nand2_1
XFILLER_202_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14523_ _07242_ _07240_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__and2_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18291_ _10248_ _09977_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__nor2_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ rbzero.debug_overlay.playerX\[0\] _04459_ _04460_ rbzero.debug_overlay.playerX\[-2\]
+ _04042_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__a221o_1
XFILLER_186_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17242_ _09812_ _09815_ _09816_ _09817_ _09819_ vssd1 vssd1 vccd1 vccd1 _09820_ sky130_fd_sc_hd__o311a_1
X_14454_ _07187_ _07190_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__and2_1
X_11666_ _04435_ _04437_ _04439_ _04440_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__o41a_1
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20356__365 clknet_1_1__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__inv_2
XFILLER_128_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13405_ _06138_ _06141_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__xor2_1
XFILLER_31_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10617_ rbzero.tex_g1\[47\] rbzero.tex_g1\[48\] _03647_ vssd1 vssd1 vccd1 vccd1 _03648_
+ sky130_fd_sc_hd__mux2_1
X_17173_ rbzero.traced_texa\[2\] _09768_ _09769_ rbzero.wall_tracer.visualWallDist\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__a22o_1
X_14385_ _06724_ _06708_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__or2_1
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ rbzero.tex_r1\[61\] rbzero.tex_r1\[60\] _04338_ vssd1 vssd1 vccd1 vccd1 _04376_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16124_ _07980_ _08102_ _08103_ vssd1 vssd1 vccd1 vccd1 _08769_ sky130_fd_sc_hd__or3_1
XFILLER_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13336_ _06071_ _06072_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__xnor2_1
X_10548_ rbzero.tex_r0\[16\] rbzero.tex_r0\[15\] _03602_ vssd1 vssd1 vccd1 vccd1 _03611_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16055_ _08679_ _08699_ vssd1 vssd1 vccd1 vccd1 _08700_ sky130_fd_sc_hd__xnor2_2
X_13267_ _05983_ _05981_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__or3_1
X_10479_ rbzero.tex_r0\[49\] rbzero.tex_r0\[48\] _03569_ vssd1 vssd1 vccd1 vccd1 _03575_
+ sky130_fd_sc_hd__mux2_1
XFILLER_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15006_ _07673_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12218_ _04886_ _04887_ _04961_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__mux2_1
XFILLER_194_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13198_ _05778_ _05934_ _05928_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__o21a_1
XFILLER_116_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19814_ rbzero.pov.ready _02821_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__and2_1
X_12149_ net50 _04907_ _04910_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__a31o_1
XFILLER_97_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03314_ clknet_0__03314_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03314_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19745_ _03100_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__clkbuf_1
X_16957_ rbzero.debug_overlay.playerY\[-2\] rbzero.debug_overlay.playerX\[-2\] _07895_
+ vssd1 vssd1 vccd1 vccd1 _09598_ sky130_fd_sc_hd__mux2_1
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15908_ _07988_ _07938_ _07939_ vssd1 vssd1 vccd1 vccd1 _08553_ sky130_fd_sc_hd__or3_1
X_19676_ _03064_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__clkbuf_1
X_16888_ _08204_ _08570_ vssd1 vssd1 vccd1 vccd1 _09529_ sky130_fd_sc_hd__nor2_1
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18627_ _02291_ _02300_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__or2b_1
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15839_ _08480_ _08481_ _08483_ vssd1 vssd1 vccd1 vccd1 _08484_ sky130_fd_sc_hd__a21bo_1
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18558_ _10239_ _09481_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__nor2_1
XFILLER_178_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17509_ _09522_ _08151_ _10074_ vssd1 vssd1 vccd1 vccd1 _10075_ sky130_fd_sc_hd__or3_1
XFILLER_166_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18489_ _01860_ _09141_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__or4_1
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 _07988_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20520_ _03413_ _03414_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__xnor2_1
XFILLER_127_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_24 rbzero.wall_tracer.visualWallDist\[-12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_46 _07939_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 net27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20451_ rbzero.texV\[-6\] _03175_ _03332_ _03356_ vssd1 vssd1 vccd1 vccd1 _01390_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_68 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20382_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__buf_1
XFILLER_107_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21003_ clknet_leaf_10_i_clk _00772_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20383__9 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__inv_2
XFILLER_130_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _04263_ vssd1 vssd1 vccd1 vccd1 _04300_
+ sky130_fd_sc_hd__mux2_1
X_20718_ clknet_leaf_62_i_clk _00008_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_157_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ _04223_ _04227_ _04228_ _04219_ _04230_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__o221a_1
XFILLER_183_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20649_ clknet_leaf_49_i_clk _00433_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10402_ _03532_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14170_ _06905_ _06906_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__nor2_1
X_11382_ rbzero.row_render.size\[3\] vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__inv_2
XFILLER_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13121_ _05761_ _05762_ _05796_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__mux2_1
X_10333_ _03496_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13052_ _05694_ _05771_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__nand2_1
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12003_ _04774_ _04777_ _04332_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__mux2_1
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17860_ _01461_ _01470_ _01468_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__a21o_1
XFILLER_79_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16811_ _09321_ _09323_ _09452_ vssd1 vssd1 vccd1 vccd1 _09453_ sky130_fd_sc_hd__o21a_1
XFILLER_121_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17791_ _10258_ _10262_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__and2_1
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19530_ _04034_ _03006_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__or2_1
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16742_ _09269_ _09273_ vssd1 vssd1 vccd1 vccd1 _09384_ sky130_fd_sc_hd__or2_1
X_13954_ _06689_ _06690_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__or2_1
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12905_ _05609_ _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__xor2_2
X_16673_ _09311_ _09312_ _09314_ vssd1 vssd1 vccd1 vccd1 _09316_ sky130_fd_sc_hd__a21oi_1
X_19461_ _02916_ _02929_ _02930_ _02911_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__o2bb2a_1
X_13885_ _05978_ _06067_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__or2_1
XFILLER_35_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18412_ _02109_ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__or2_1
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ rbzero.wall_tracer.visualWallDist\[9\] _05571_ _05572_ vssd1 vssd1 vccd1
+ vccd1 _05573_ sky130_fd_sc_hd__a21o_1
X_15624_ rbzero.wall_tracer.stepDistX\[-1\] vssd1 vssd1 vccd1 vccd1 _08269_ sky130_fd_sc_hd__inv_2
X_19392_ _02868_ _02871_ _02869_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a21bo_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18343_ _09141_ _01620_ _02041_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__or3_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ rbzero.wall_tracer.stepDistY\[0\] vssd1 vssd1 vccd1 vccd1 _08200_ sky130_fd_sc_hd__inv_2
XFILLER_187_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12767_ rbzero.map_rom.f1 _05512_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__or2_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14506_ _07237_ _07240_ _07242_ vssd1 vssd1 vccd1 vccd1 _07243_ sky130_fd_sc_hd__a21boi_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18274_ _01646_ _01883_ _10271_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__a21oi_1
X_11718_ _04480_ _04490_ _04492_ _04496_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__o22a_1
X_15486_ _08127_ _08130_ vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__nor2_1
XFILLER_159_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ _05416_ _05442_ _05443_ _05444_ _05445_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__a311o_1
XFILLER_202_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14437_ _07110_ _07173_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__xnor2_1
X_17225_ _08937_ _09803_ vssd1 vssd1 vccd1 vccd1 _09804_ sky130_fd_sc_hd__xor2_1
XFILLER_128_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput11 i_gpout1_sel[3] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__buf_8
X_11649_ _04422_ _04427_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nor2_1
Xinput22 i_gpout3_sel[2] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_6
XFILLER_156_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput33 i_gpout5_sel[1] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_4
XFILLER_168_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput44 i_reset_lock_a vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__buf_6
X_17156_ _07679_ vssd1 vssd1 vccd1 vccd1 _09767_ sky130_fd_sc_hd__clkbuf_4
XFILLER_196_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14368_ _07104_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__inv_2
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16107_ _08743_ _08750_ _08751_ vssd1 vssd1 vccd1 vccd1 _08752_ sky130_fd_sc_hd__a21oi_1
X_13319_ _05922_ _06054_ _06055_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__a21o_1
X_17087_ _09579_ _09581_ vssd1 vssd1 vccd1 vccd1 _09727_ sky130_fd_sc_hd__and2b_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14299_ _06842_ _06881_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__xor2_1
XFILLER_157_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16038_ _08680_ _08681_ vssd1 vssd1 vccd1 vccd1 _08683_ sky130_fd_sc_hd__xnor2_1
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17989_ _01688_ _01690_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__nand2_1
XFILLER_81_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19728_ _03091_ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_26_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19659_ _03055_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__clkbuf_1
XFILLER_93_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21621_ clknet_leaf_73_i_clk _01390_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-6\] sky130_fd_sc_hd__dfxtp_1
X_21552_ net473 _01321_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20503_ _09750_ _03399_ _03400_ _03250_ rbzero.texV\[2\] vssd1 vssd1 vccd1 vccd1
+ _01398_ sky130_fd_sc_hd__a32o_1
XFILLER_119_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21483_ net404 _01252_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20434_ rbzero.texV\[-9\] _03175_ _03332_ _03342_ vssd1 vssd1 vccd1 vccd1 _01387_
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10951_ rbzero.tex_b1\[16\] rbzero.tex_b1\[17\] _03817_ vssd1 vssd1 vccd1 vccd1 _03823_
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13670_ _06406_ _06078_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__or2_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10882_ rbzero.tex_b1\[49\] rbzero.tex_b1\[50\] _03784_ vssd1 vssd1 vccd1 vccd1 _03787_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ rbzero.map_rom.c6 _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__and2_1
XFILLER_25_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15340_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07985_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _05304_ _05305_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__nor2_1
XFILLER_8_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11503_ rbzero.tex_r0\[7\] rbzero.tex_r0\[6\] _04273_ vssd1 vssd1 vccd1 vccd1 _04283_
+ sky130_fd_sc_hd__mux2_1
X_15271_ _05495_ _07914_ _07915_ _05195_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__o211a_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12483_ rbzero.wall_tracer.trackDistX\[-7\] vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__03317_ clknet_0__03317_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03317_
+ sky130_fd_sc_hd__clkbuf_16
X_17010_ _09647_ _09649_ vssd1 vssd1 vccd1 vccd1 _09650_ sky130_fd_sc_hd__nor2_1
X_14222_ _06955_ _06957_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__nand2_1
XFILLER_172_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11434_ _04213_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__clkbuf_4
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14153_ _06741_ _06888_ _06889_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__a21bo_1
X_11365_ _04141_ _04142_ _04143_ _04144_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__or4_1
X_13104_ _05634_ _05636_ _05796_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__mux2_1
X_10316_ _03487_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__clkbuf_1
X_14084_ _06799_ _06814_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__xnor2_1
X_18961_ _02610_ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11296_ _04073_ _04072_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__nand2_1
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17912_ _01516_ _01522_ _01614_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__a21oi_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _05760_ _05763_ _05767_ _05769_ _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__o2111ai_2
XFILLER_152_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18892_ _02561_ rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_cmd\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__or3b_1
XFILLER_117_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17843_ _01442_ _01546_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17774_ _08202_ _01476_ _08417_ _08445_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14986_ _00008_ _07552_ _07663_ vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__a21oi_1
X_19513_ _02973_ _02979_ _02989_ _03913_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__a31o_1
X_16725_ _09365_ _09366_ vssd1 vssd1 vccd1 vccd1 _09367_ sky130_fd_sc_hd__nand2_1
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13937_ _06161_ _06667_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__nor2_2
XFILLER_207_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19444_ rbzero.debug_overlay.vplaneY\[-1\] rbzero.debug_overlay.vplaneY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__or2_1
X_16656_ _09282_ _09297_ _09298_ vssd1 vssd1 vccd1 vccd1 _09299_ sky130_fd_sc_hd__nand3_1
X_13868_ _06604_ _06554_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_0__03044_ _03044_ vssd1 vssd1 vccd1 vccd1 clknet_0__03044_ sky130_fd_sc_hd__clkbuf_16
X_15607_ _08245_ _08251_ vssd1 vssd1 vccd1 vccd1 _08252_ sky130_fd_sc_hd__xor2_1
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12819_ rbzero.wall_tracer.mapY\[10\] _05404_ _05555_ vssd1 vssd1 vccd1 vccd1 _05557_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_50_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19375_ _02851_ _02855_ _02852_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__o21ai_1
X_16587_ _09224_ _09229_ vssd1 vssd1 vccd1 vccd1 _09230_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13799_ _06057_ _06061_ vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__nor2_1
XFILLER_72_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18326_ _01905_ _02013_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__or2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15538_ _08181_ _08182_ _07970_ vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__a21o_1
XFILLER_124_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18257_ _01498_ _08423_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__nor2_1
X_15469_ _08111_ _08022_ _08113_ vssd1 vssd1 vccd1 vccd1 _08114_ sky130_fd_sc_hd__o21ai_1
XFILLER_124_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17208_ _09779_ _09789_ _09790_ _09781_ rbzero.wall_tracer.mapX\[8\] vssd1 vssd1
+ vccd1 vccd1 _00573_ sky130_fd_sc_hd__a32o_1
XFILLER_200_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18188_ _01753_ _01769_ _01768_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a21bo_1
XFILLER_128_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _07530_ _09763_ rbzero.row_render.size\[2\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00530_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20983_ clknet_leaf_10_i_clk _00752_ vssd1 vssd1 vccd1 vccd1 rbzero.color_floor\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21604_ net145 _01373_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[55\] sky130_fd_sc_hd__dfxtp_1
XFILLER_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21535_ net456 _01304_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21466_ net387 _01235_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20417_ rbzero.traced_texa\[-11\] rbzero.texV\[-11\] vssd1 vssd1 vccd1 vccd1 _03328_
+ sky130_fd_sc_hd__or2_1
XFILLER_181_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21397_ net318 _01166_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11150_ _03923_ _03928_ _03932_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__or4_2
XFILLER_190_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11081_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _03887_ vssd1 vssd1 vccd1 vccd1 _03891_
+ sky130_fd_sc_hd__mux2_1
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ rbzero.wall_tracer.stepDistY\[2\] _07562_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07563_ sky130_fd_sc_hd__mux2_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14771_ _05844_ _05952_ _07469_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__and3_1
X_11983_ _04755_ _04756_ _04757_ _04247_ _04332_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__o221a_1
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16510_ _08995_ _08997_ vssd1 vssd1 vccd1 vccd1 _09154_ sky130_fd_sc_hd__nor2_1
X_13722_ _06427_ _06457_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10934_ rbzero.tex_b1\[24\] rbzero.tex_b1\[25\] _03806_ vssd1 vssd1 vccd1 vccd1 _03814_
+ sky130_fd_sc_hd__mux2_1
X_17490_ _08335_ _09703_ vssd1 vssd1 vccd1 vccd1 _10056_ sky130_fd_sc_hd__and2_1
XFILLER_186_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16441_ rbzero.wall_tracer.texu\[0\] _09085_ vssd1 vssd1 vccd1 vccd1 _09086_ sky130_fd_sc_hd__or2_1
X_13653_ _06283_ _06389_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__and2_1
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ rbzero.tex_b1\[57\] rbzero.tex_b1\[58\] _03773_ vssd1 vssd1 vccd1 vccd1 _03778_
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _05289_ _05357_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__nand2_1
X_16372_ _09013_ _09015_ vssd1 vssd1 vccd1 vccd1 _09017_ sky130_fd_sc_hd__and2_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19160_ _05189_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__buf_6
XFILLER_13_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13584_ _06308_ _06320_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__xnor2_2
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _03740_ vssd1 vssd1 vccd1 vccd1 _03742_
+ sky130_fd_sc_hd__mux2_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _01807_ _01810_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__or2_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _07959_ _07967_ vssd1 vssd1 vccd1 vccd1 _07968_ sky130_fd_sc_hd__nor2_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12535_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__or2_2
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19091_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.spi_buffer\[0\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__mux2_1
XFILLER_173_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18042_ _09668_ _09693_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__nor2_1
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15254_ rbzero.debug_overlay.playerX\[-6\] _07897_ vssd1 vssd1 vccd1 vccd1 _07899_
+ sky130_fd_sc_hd__nand2_1
X_12466_ rbzero.wall_tracer.trackDistY\[7\] _05218_ _05220_ rbzero.wall_tracer.trackDistX\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14205_ _06664_ _06940_ _06941_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__a21oi_1
X_11417_ _04022_ _04187_ _04186_ gpout0.hpos\[5\] _04196_ vssd1 vssd1 vccd1 vccd1
+ _04197_ sky130_fd_sc_hd__o221a_1
X_15185_ _07837_ _07838_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__xnor2_1
X_12397_ _05157_ _05160_ _05163_ net34 net35 vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__a32o_1
XFILLER_67_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14136_ _06861_ _06871_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__nand2_1
X_11348_ _04088_ _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__nand2_1
XFILLER_119_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19993_ rbzero.pov.ready_buffer\[19\] _03252_ _03253_ _07730_ _03254_ vssd1 vssd1
+ vccd1 vccd1 _01034_ sky130_fd_sc_hd__o221a_1
XFILLER_67_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14067_ _06769_ _06707_ vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__or2_1
X_18944_ _02601_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11279_ _04057_ _04058_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__nand2_1
X_13018_ _05743_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__or2_1
XFILLER_140_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18875_ _02546_ _02547_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17826_ _01523_ _01529_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17757_ _01459_ _01460_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14969_ _07654_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16708_ rbzero.wall_tracer.visualWallDist\[9\] _04015_ vssd1 vssd1 vccd1 vccd1 _09350_
+ sky130_fd_sc_hd__nand2_4
XFILLER_35_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17688_ _10236_ _10252_ vssd1 vssd1 vccd1 vccd1 _10253_ sky130_fd_sc_hd__xor2_2
XFILLER_207_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19427_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.debug_overlay.vplaneY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__nor2_1
X_16639_ _09277_ _09281_ vssd1 vssd1 vccd1 vccd1 _09282_ sky130_fd_sc_hd__xor2_1
XFILLER_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20221__243 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__inv_2
XFILLER_167_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19358_ _07703_ _02846_ _02847_ _07706_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__a31o_1
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18309_ _02006_ _02008_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__xnor2_1
XFILLER_200_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19289_ rbzero.spi_registers.got_new_leak _02730_ _02728_ _02799_ vssd1 vssd1 vccd1
+ vccd1 _00785_ sky130_fd_sc_hd__a31o_1
XFILLER_136_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21320_ net241 _01089_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21251_ clknet_leaf_91_i_clk _01020_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_85_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21182_ clknet_leaf_7_i_clk _00951_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20304__318 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__inv_2
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20966_ clknet_leaf_8_i_clk _00735_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_26_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20897_ clknet_leaf_68_i_clk _00666_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10650_ rbzero.tex_g1\[31\] rbzero.tex_g1\[32\] _03658_ vssd1 vssd1 vccd1 vccd1 _03665_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20196__220 clknet_1_1__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__inv_2
XFILLER_10_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10581_ _03628_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12320_ _05087_ _04666_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__nand2_1
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21518_ net439 _01287_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ _04325_ _04965_ _04976_ _05020_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__o2bb2a_2
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21449_ net370 _01218_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11202_ _03924_ _03925_ rbzero.map_rom.a6 rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1
+ _03991_ sky130_fd_sc_hd__o22a_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12182_ _04948_ _04952_ net12 vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__o21ai_1
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11133_ rbzero.debug_overlay.playerX\[0\] _03919_ _03921_ rbzero.debug_overlay.playerY\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__a2bb2o_1
X_16990_ _09628_ _09629_ vssd1 vssd1 vccd1 vccd1 _09630_ sky130_fd_sc_hd__and2b_1
XFILLER_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15941_ _08535_ _08536_ vssd1 vssd1 vccd1 vccd1 _08586_ sky130_fd_sc_hd__xnor2_1
XFILLER_62_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11064_ rbzero.tex_b0\[27\] rbzero.tex_b0\[26\] _03876_ vssd1 vssd1 vccd1 vccd1 _03882_
+ sky130_fd_sc_hd__mux2_1
XFILLER_114_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18660_ _01498_ _01860_ _09027_ _09350_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__or4_1
XFILLER_76_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15872_ _08448_ _08516_ vssd1 vssd1 vccd1 vccd1 _08517_ sky130_fd_sc_hd__xor2_2
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17611_ _10031_ _10033_ _10174_ _10175_ vssd1 vssd1 vccd1 vccd1 _10177_ sky130_fd_sc_hd__o211ai_2
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14823_ rbzero.wall_tracer.stepDistY\[-2\] _07461_ vssd1 vssd1 vccd1 vccd1 _07550_
+ sky130_fd_sc_hd__nor2_1
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18591_ _02250_ _02287_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__xor2_1
XFILLER_64_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17542_ _10092_ _10107_ vssd1 vssd1 vccd1 vccd1 _10108_ sky130_fd_sc_hd__xor2_2
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14754_ _05794_ _07104_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__nor2_1
XFILLER_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11966_ _04739_ _04740_ _04329_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__mux2_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13705_ _06402_ _06403_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10917_ rbzero.tex_b1\[32\] rbzero.tex_b1\[33\] _03795_ vssd1 vssd1 vccd1 vccd1 _03805_
+ sky130_fd_sc_hd__mux2_1
X_17473_ _09908_ _09917_ _09915_ vssd1 vssd1 vccd1 vccd1 _10039_ sky130_fd_sc_hd__a21o_1
X_14685_ _07394_ _07421_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__nand2_1
X_11897_ rbzero.tex_b0\[10\] _04213_ _04329_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__a21o_1
XFILLER_44_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19212_ rbzero.color_floor\[1\] _02751_ _02754_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__a21o_1
XFILLER_60_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13636_ _06349_ _06372_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__xnor2_2
XFILLER_73_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16424_ _08951_ _08953_ vssd1 vssd1 vccd1 vccd1 _09069_ sky130_fd_sc_hd__xor2_4
XFILLER_177_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10848_ rbzero.tex_g0\[2\] rbzero.tex_g0\[1\] _03762_ vssd1 vssd1 vccd1 vccd1 _03769_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19143_ _02709_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__buf_2
X_16355_ _08358_ _08365_ _08999_ vssd1 vssd1 vccd1 vccd1 _09000_ sky130_fd_sc_hd__a21o_2
X_13567_ _06111_ _06128_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__xnor2_2
X_10779_ rbzero.tex_g0\[35\] rbzero.tex_g0\[34\] _03729_ vssd1 vssd1 vccd1 vccd1 _03733_
+ sky130_fd_sc_hd__mux2_1
XFILLER_118_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15306_ _07904_ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__buf_4
X_12518_ _05272_ _05253_ _05261_ _05262_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__a211o_1
X_16286_ _08909_ _08853_ vssd1 vssd1 vccd1 vccd1 _08931_ sky130_fd_sc_hd__or2b_1
X_19074_ _02669_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__clkbuf_1
X_13498_ _06168_ _06208_ _06234_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__a21o_1
XFILLER_195_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18025_ _01724_ _01725_ _01716_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__o21ai_1
X_12449_ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__buf_8
X_15237_ _07881_ _07868_ _07872_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__and3b_1
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15168_ _07818_ _07819_ _07822_ vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__and3_1
XFILLER_114_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _06855_ _06699_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__and2b_1
XFILLER_99_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19976_ rbzero.pov.ready_buffer\[27\] _03240_ _03243_ rbzero.debug_overlay.facingY\[-4\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__o221a_1
X_15099_ rbzero.debug_overlay.vplaneX\[10\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__nand2_1
XFILLER_87_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18927_ _02591_ vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18858_ _02530_ _02531_ _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17809_ _01494_ _01512_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__xor2_2
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18789_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.stepDistY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__and2_1
X_20820_ clknet_leaf_49_i_clk _00589_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20751_ clknet_leaf_38_i_clk _00520_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_63_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20682_ clknet_leaf_50_i_clk _00466_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_50_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21303_ net224 _01072_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21234_ clknet_leaf_18_i_clk _01003_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21165_ clknet_leaf_89_i_clk _00934_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20116_ clknet_1_1__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__buf_1
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21096_ net186 _00865_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20047_ _04990_ _04322_ _03275_ _03911_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__a31o_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20228__249 clknet_1_0__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__inv_2
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _04595_ _04596_ _04345_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__mux2_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ rbzero.tex_g0\[10\] _04212_ _04217_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__a21o_1
XFILLER_121_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20949_ clknet_leaf_2_i_clk _00718_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_cmd\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10702_ _03692_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14470_ _07131_ _07205_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__and2_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ rbzero.debug_overlay.vplaneX\[0\] _04459_ _04460_ rbzero.debug_overlay.vplaneX\[-2\]
+ gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__a221o_1
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13421_ _06002_ _05976_ _06004_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__a21bo_1
X_10633_ rbzero.tex_g1\[39\] rbzero.tex_g1\[40\] _03647_ vssd1 vssd1 vccd1 vccd1 _03656_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16140_ _08674_ _08112_ _08747_ vssd1 vssd1 vccd1 vccd1 _08785_ sky130_fd_sc_hd__or3_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13352_ _06077_ _06088_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10564_ _03619_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_154_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12303_ net23 net22 _05071_ net24 vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__a31o_1
X_16071_ _08696_ _08714_ vssd1 vssd1 vccd1 vccd1 _08716_ sky130_fd_sc_hd__nor2_1
XFILLER_155_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13283_ _06006_ _06019_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__xnor2_1
X_10495_ _03583_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__clkbuf_1
X_15022_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__nand2_1
X_12234_ net17 net16 _05003_ net18 vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a31o_1
X_19830_ rbzero.pov.ready_buffer\[61\] _07999_ _03146_ vssd1 vssd1 vccd1 vccd1 _03150_
+ sky130_fd_sc_hd__mux2_1
X_12165_ net48 _04903_ _04922_ net40 _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a221o_1
XFILLER_190_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11116_ rbzero.tex_b0\[2\] rbzero.tex_b0\[1\] _03557_ vssd1 vssd1 vccd1 vccd1 _03909_
+ sky130_fd_sc_hd__mux2_1
XFILLER_116_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19761_ rbzero.pov.spi_buffer\[54\] rbzero.pov.spi_buffer\[55\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03109_ sky130_fd_sc_hd__mux2_1
X_12096_ _04867_ _04837_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__and2_1
X_16973_ _09609_ _09612_ vssd1 vssd1 vccd1 vccd1 _09613_ sky130_fd_sc_hd__xnor2_2
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18712_ _02398_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__buf_4
XFILLER_110_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15924_ _08497_ _08501_ vssd1 vssd1 vccd1 vccd1 _08569_ sky130_fd_sc_hd__xnor2_2
X_11047_ rbzero.tex_b0\[35\] rbzero.tex_b0\[34\] _03865_ vssd1 vssd1 vccd1 vccd1 _03873_
+ sky130_fd_sc_hd__mux2_1
X_19692_ rbzero.pov.spi_buffer\[21\] rbzero.pov.spi_buffer\[22\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03073_ sky130_fd_sc_hd__mux2_1
XFILLER_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 i_gpout1_sel[1] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_6
X_18643_ _08418_ _02336_ _02338_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__03292_ _03292_ vssd1 vssd1 vccd1 vccd1 clknet_0__03292_ sky130_fd_sc_hd__clkbuf_16
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _08109_ _08042_ _08125_ _08084_ vssd1 vssd1 vccd1 vccd1 _08500_ sky130_fd_sc_hd__o22ai_1
XFILLER_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _07487_ _07456_ _07533_ _07535_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__a211oi_4
XFILLER_91_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18574_ _02188_ _02190_ _02187_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a21bo_1
XFILLER_18_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15786_ _08330_ _08415_ _08429_ vssd1 vssd1 vccd1 vccd1 _08431_ sky130_fd_sc_hd__a21oi_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _05721_ _05734_ _05707_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__or3_1
XFILLER_75_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17525_ _09979_ _09984_ vssd1 vssd1 vccd1 vccd1 _10091_ sky130_fd_sc_hd__and2_1
XFILLER_51_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14737_ _05844_ _07471_ _06239_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__a21o_1
X_11949_ rbzero.tex_b0\[33\] rbzero.tex_b0\[32\] _04356_ vssd1 vssd1 vccd1 vccd1 _04725_
+ sky130_fd_sc_hd__mux2_1
XFILLER_162_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17456_ _09614_ _10022_ vssd1 vssd1 vccd1 vccd1 _10023_ sky130_fd_sc_hd__xnor2_4
XFILLER_20_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14668_ _07394_ _07399_ _07404_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__or3b_1
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16407_ _08412_ _08438_ _09051_ vssd1 vssd1 vccd1 vccd1 _09052_ sky130_fd_sc_hd__a21oi_2
XFILLER_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _05823_ _05920_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__or2_2
XFILLER_193_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17387_ _09952_ _09953_ vssd1 vssd1 vccd1 vccd1 _09954_ sky130_fd_sc_hd__nand2_1
XFILLER_125_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14599_ _07218_ _07323_ _07331_ _07216_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__a211o_1
XFILLER_186_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19126_ net41 rbzero.spi_registers.ss_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02698_ sky130_fd_sc_hd__mux2_1
XFILLER_158_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16338_ _07566_ _07568_ _07571_ _08220_ vssd1 vssd1 vccd1 vccd1 _08983_ sky130_fd_sc_hd__or4_2
XFILLER_118_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19057_ rbzero.pov.spi_buffer\[59\] rbzero.pov.ready_buffer\[59\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02661_ sky130_fd_sc_hd__mux2_1
X_16269_ _08250_ _08331_ _08862_ vssd1 vssd1 vccd1 vccd1 _08914_ sky130_fd_sc_hd__a21oi_1
X_20333__344 clknet_1_1__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__inv_2
XFILLER_145_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18008_ _01708_ _01709_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__nand2_1
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19959_ _03246_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__clkbuf_4
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20803_ clknet_leaf_30_i_clk _00572_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_150_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20734_ clknet_leaf_81_i_clk _00503_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_81_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20665_ clknet_leaf_62_i_clk _00449_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20596_ rbzero.wall_tracer.rayAddendY\[-7\] _03443_ _07756_ _03461_ vssd1 vssd1 vccd1
+ vccd1 _01430_ sky130_fd_sc_hd__a22o_1
XFILLER_109_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_96_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21217_ clknet_leaf_20_i_clk _00986_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21148_ clknet_leaf_87_i_clk _00917_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_20058__96 clknet_1_1__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__inv_2
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13970_ _06614_ _06706_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__nand2_2
X_21079_ net169 _00848_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _05567_ _05576_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__nor2_1
XFILLER_132_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_34_i_clk clknet_opt_6_1_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15640_ _08282_ _08283_ _08284_ _07996_ vssd1 vssd1 vccd1 vccd1 _08285_ sky130_fd_sc_hd__o22ai_1
XFILLER_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ rbzero.wall_tracer.rayAddendX\[-2\] _05588_ _05560_ vssd1 vssd1 vccd1 vccd1
+ _05589_ sky130_fd_sc_hd__mux2_2
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19620__73 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__inv_2
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ rbzero.tex_g0\[33\] rbzero.tex_g0\[32\] _04341_ vssd1 vssd1 vccd1 vccd1 _04581_
+ sky130_fd_sc_hd__mux2_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _08214_ _08215_ vssd1 vssd1 vccd1 vccd1 _08216_ sky130_fd_sc_hd__nor2_2
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _05513_ _05519_ _05520_ _05512_ rbzero.map_rom.i_col\[4\] vssd1 vssd1 vccd1
+ vccd1 _05527_ sky130_fd_sc_hd__a32o_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ rbzero.wall_tracer.trackDistX\[-3\] rbzero.wall_tracer.stepDistX\[-3\] vssd1
+ vssd1 vccd1 vccd1 _09880_ sky130_fd_sc_hd__or2_1
XFILLER_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14522_ _07258_ _07053_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__xnor2_1
X_11734_ rbzero.debug_overlay.playerX\[-8\] _04466_ _04499_ rbzero.debug_overlay.playerX\[4\]
+ _04512_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__a221o_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _01988_ _01989_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__xnor2_1
XFILLER_30_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_49_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17241_ _08940_ _08943_ _09818_ vssd1 vssd1 vccd1 vccd1 _09819_ sky130_fd_sc_hd__o21ai_1
XFILLER_202_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11665_ gpout0.hpos\[8\] _04443_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__and2_2
X_14453_ _07188_ _07189_ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__and2b_1
XFILLER_70_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10616_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__clkbuf_4
X_13404_ _06139_ _06140_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__xnor2_1
X_14384_ _06696_ _06740_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__or2_1
X_17172_ rbzero.traced_texa\[1\] _09768_ _09769_ rbzero.wall_tracer.visualWallDist\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a22o_1
X_11596_ rbzero.tex_r1\[63\] rbzero.tex_r1\[62\] _04338_ vssd1 vssd1 vccd1 vccd1 _04375_
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16123_ _08008_ _08128_ vssd1 vssd1 vccd1 vccd1 _08768_ sky130_fd_sc_hd__or2_1
X_13335_ _06059_ _06060_ _06045_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__a21oi_1
X_10547_ _03610_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266_ _06002_ _05976_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__xnor2_1
X_16054_ _08676_ _08677_ vssd1 vssd1 vccd1 vccd1 _08699_ sky130_fd_sc_hd__xor2_1
X_10478_ _03574_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12217_ _04883_ _04884_ _04966_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__mux2_1
X_15005_ rbzero.wall_tracer.stepDistX\[9\] _07582_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07673_ sky130_fd_sc_hd__mux2_1
XFILLER_170_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13197_ _05867_ _05688_ _05801_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__mux2_1
XFILLER_68_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19813_ _03135_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__clkbuf_1
X_12148_ net49 _04903_ _04918_ net52 vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__a22o_1
XFILLER_123_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03313_ clknet_0__03313_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03313_
+ sky130_fd_sc_hd__clkbuf_16
X_19744_ rbzero.pov.spi_buffer\[46\] rbzero.pov.spi_buffer\[47\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03100_ sky130_fd_sc_hd__mux2_1
X_12079_ net5 _04850_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__nor2_1
X_16956_ _09594_ _09596_ vssd1 vssd1 vccd1 vccd1 _09597_ sky130_fd_sc_hd__xor2_4
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15907_ _08551_ _08481_ vssd1 vssd1 vccd1 vccd1 _08552_ sky130_fd_sc_hd__xor2_1
X_19675_ rbzero.pov.spi_buffer\[13\] rbzero.pov.spi_buffer\[14\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03064_ sky130_fd_sc_hd__mux2_1
X_16887_ _09525_ _09527_ vssd1 vssd1 vccd1 vccd1 _09528_ sky130_fd_sc_hd__and2_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18626_ _02316_ _02322_ rbzero.wall_tracer.trackDistX\[10\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00599_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _07923_ _07967_ _08482_ vssd1 vssd1 vccd1 vccd1 _08483_ sky130_fd_sc_hd__or3_1
XFILLER_53_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18557_ _02144_ _02158_ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__a21bo_1
X_15769_ _08408_ _08402_ vssd1 vssd1 vccd1 vccd1 _08414_ sky130_fd_sc_hd__or2b_1
XFILLER_45_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17508_ _07974_ _08158_ vssd1 vssd1 vccd1 vccd1 _10074_ sky130_fd_sc_hd__or2_1
XFILLER_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18488_ _02039_ _02042_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__nand2_1
XFILLER_162_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17439_ _10003_ _10005_ vssd1 vssd1 vccd1 vccd1 _10006_ sky130_fd_sc_hd__xnor2_2
XANTENNA_14 _08037_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_25 rbzero.wall_tracer.visualWallDist\[-7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _08096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_58 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20450_ _03353_ _03355_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__xnor2_1
XANTENNA_69 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19109_ rbzero.spi_registers.spi_buffer\[10\] rbzero.spi_registers.spi_buffer\[9\]
+ _02676_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__mux2_1
XFILLER_192_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21002_ clknet_leaf_8_i_clk _00771_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_sky
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20717_ clknet_leaf_46_i_clk _00007_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11450_ _04229_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__buf_4
X_20648_ clknet_leaf_57_i_clk _00432_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ rbzero.tex_r1\[19\] rbzero.tex_r1\[20\] _03527_ vssd1 vssd1 vccd1 vccd1 _03532_
+ sky130_fd_sc_hd__mux2_1
X_11381_ rbzero.row_render.size\[4\] vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__inv_2
X_20579_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__or2_1
XFILLER_180_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13120_ _05690_ _05801_ _05817_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__o21ai_1
XFILLER_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10332_ rbzero.tex_r1\[52\] rbzero.tex_r1\[53\] _03494_ vssd1 vssd1 vccd1 vccd1 _03496_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _05780_ _05746_ _05782_ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__nand4_2
XFILLER_133_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12002_ _04775_ _04776_ _04218_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__mux2_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16810_ _09318_ _09320_ vssd1 vssd1 vccd1 vccd1 _09452_ sky130_fd_sc_hd__or2_1
XFILLER_87_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17790_ _10243_ _10251_ _01493_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__a21o_1
XFILLER_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16741_ _09251_ _09261_ _09259_ vssd1 vssd1 vccd1 vccd1 _09383_ sky130_fd_sc_hd__a21o_1
XFILLER_120_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13953_ _06610_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__clkbuf_4
XFILLER_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19460_ _02940_ _02941_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__nor2_1
X_12904_ _05562_ _05566_ _05619_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__and3_1
X_20362__370 clknet_1_0__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__inv_2
X_16672_ _09311_ _09312_ _09314_ vssd1 vssd1 vccd1 vccd1 _09315_ sky130_fd_sc_hd__and3_1
X_13884_ _06201_ _06052_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__nor2_1
XFILLER_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18411_ _01946_ _01949_ _02108_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__and3_1
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15623_ _08191_ _08265_ _08267_ vssd1 vssd1 vccd1 vccd1 _08268_ sky130_fd_sc_hd__a21bo_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ _07728_ _02872_ _02877_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__a21o_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _04031_ _05327_ _05371_ _04001_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__a31o_1
XFILLER_188_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _02039_ _02040_ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__nand2_1
XFILLER_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _08196_ _08198_ _07951_ vssd1 vssd1 vccd1 vccd1 _08199_ sky130_fd_sc_hd__a21o_2
XFILLER_199_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _05496_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__buf_2
XFILLER_203_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14505_ _07238_ _07241_ _07239_ _07075_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__a22o_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _01646_ _01972_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11717_ rbzero.debug_overlay.facingX\[10\] _04453_ _04493_ _04495_ vssd1 vssd1 vccd1
+ vccd1 _04496_ sky130_fd_sc_hd__a211o_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15485_ _08047_ _08124_ _08128_ _08129_ vssd1 vssd1 vccd1 vccd1 _08130_ sky130_fd_sc_hd__o22a_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12697_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] vssd1
+ vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__xnor2_2
XFILLER_188_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17224_ _08939_ _08851_ vssd1 vssd1 vccd1 vccd1 _09803_ sky130_fd_sc_hd__and2_1
XFILLER_35_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14436_ _06689_ _06760_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__nor2_1
X_11648_ gpout0.hpos\[5\] _04424_ _04426_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__or3_1
XFILLER_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 i_gpout1_sel[4] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_6
XFILLER_35_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput23 i_gpout3_sel[3] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_6
Xinput34 i_gpout5_sel[2] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_6
XFILLER_196_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17155_ rbzero.row_render.texu\[5\] _09766_ _07728_ rbzero.wall_tracer.texu\[5\]
+ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__a22o_1
Xinput45 i_reset_lock_b vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_6
X_11579_ rbzero.tex_r1\[17\] rbzero.tex_r1\[16\] _04290_ vssd1 vssd1 vccd1 vccd1 _04358_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14367_ _05779_ _07103_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__or2_2
XFILLER_7_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16106_ _08744_ _08749_ vssd1 vssd1 vccd1 vccd1 _08751_ sky130_fd_sc_hd__nor2_1
XFILLER_157_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13318_ _05973_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__inv_2
X_17086_ _09657_ _09725_ vssd1 vssd1 vccd1 vccd1 _09726_ sky130_fd_sc_hd__xnor2_2
X_14298_ _06882_ _07034_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__and2_1
XFILLER_196_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16037_ _08680_ _08681_ vssd1 vssd1 vccd1 vccd1 _08682_ sky130_fd_sc_hd__or2_1
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13249_ _05962_ _05976_ _05985_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__a21o_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17988_ _01689_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__inv_2
XFILLER_57_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19727_ rbzero.pov.spi_buffer\[38\] rbzero.pov.spi_buffer\[39\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03091_ sky130_fd_sc_hd__mux2_1
X_16939_ _09442_ _09443_ vssd1 vssd1 vccd1 vccd1 _09580_ sky130_fd_sc_hd__nor2_1
XFILLER_133_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19658_ rbzero.pov.spi_buffer\[5\] rbzero.pov.spi_buffer\[6\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
XFILLER_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18609_ _02109_ _02213_ _02211_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__a21oi_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21620_ clknet_leaf_73_i_clk _01389_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21551_ net472 _01320_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20502_ _03395_ _03396_ _03397_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__a21o_1
X_21482_ net403 _01251_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20433_ _03340_ _03341_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20190__215 clknet_1_0__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__inv_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10950_ _03822_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_95_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10881_ _03786_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12620_ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__clkbuf_4
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__and2_1
XFILLER_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11502_ rbzero.tex_r0\[5\] rbzero.tex_r0\[4\] _04273_ vssd1 vssd1 vccd1 vccd1 _04282_
+ sky130_fd_sc_hd__mux2_1
XFILLER_145_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15270_ rbzero.debug_overlay.playerX\[-5\] _05495_ vssd1 vssd1 vccd1 vccd1 _07915_
+ sky130_fd_sc_hd__nand2_1
X_12482_ rbzero.wall_tracer.trackDistX\[-6\] vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__03316_ clknet_0__03316_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03316_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11433_ _04212_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__buf_4
X_14221_ _06955_ _06957_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__nor2_1
XFILLER_165_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152_ _05825_ _06740_ _06678_ _06704_ vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__o22ai_1
XFILLER_165_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11364_ _03476_ _04025_ gpout0.hpos\[9\] vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__o21ba_4
XFILLER_138_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10315_ rbzero.tex_r1\[60\] rbzero.tex_r1\[61\] _03483_ vssd1 vssd1 vccd1 vccd1 _03487_
+ sky130_fd_sc_hd__mux2_1
X_13103_ _05838_ _05839_ _05811_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__mux2_1
X_14083_ _06703_ _06819_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__nor2_1
X_18960_ rbzero.pov.spi_buffer\[13\] rbzero.pov.ready_buffer\[13\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02610_ sky130_fd_sc_hd__mux2_1
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11295_ _04071_ _04074_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__nor2_1
XFILLER_152_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17911_ _01517_ _01521_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__and2_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _05701_ _05702_ _05683_ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__or4_1
XFILLER_106_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18891_ rbzero.spi_registers.spi_cmd\[1\] rbzero.spi_registers.spi_cmd\[0\] vssd1
+ vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__or2_1
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17842_ _01543_ _01545_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17773_ _01474_ _08202_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__or4_1
XFILLER_47_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14985_ rbzero.wall_tracer.stepDistX\[-1\] _07650_ vssd1 vssd1 vccd1 vccd1 _07663_
+ sky130_fd_sc_hd__nor2_1
X_19512_ _02973_ _02979_ _02989_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a21oi_1
XFILLER_75_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16724_ _08821_ _08159_ _08151_ _09243_ vssd1 vssd1 vccd1 vccd1 _09366_ sky130_fd_sc_hd__o22ai_1
XFILLER_35_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13936_ _06245_ _06672_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__nor2_1
XFILLER_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19443_ _02923_ _02924_ _02921_ _02922_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__o211a_1
X_16655_ _09291_ _09293_ _09296_ vssd1 vssd1 vccd1 vccd1 _09298_ sky130_fd_sc_hd__a21o_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13867_ _06464_ _06552_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__nand2_1
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03043_ _03043_ vssd1 vssd1 vccd1 vccd1 clknet_0__03043_ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15606_ _08217_ _08225_ _08250_ vssd1 vssd1 vccd1 vccd1 _08251_ sky130_fd_sc_hd__o21a_1
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19374_ _02860_ _02861_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__nand2_1
X_12818_ _05533_ _05555_ _05556_ _05284_ rbzero.wall_tracer.mapY\[10\] vssd1 vssd1
+ vccd1 vccd1 _00417_ sky130_fd_sc_hd__a32o_1
X_16586_ _09227_ _09228_ vssd1 vssd1 vccd1 vccd1 _09229_ sky130_fd_sc_hd__xor2_1
XFILLER_15_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13798_ _05877_ _05888_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__nor2_1
XFILLER_203_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18325_ _01801_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__and2_1
XFILLER_163_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15537_ _07560_ _08171_ _07562_ vssd1 vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__o21ai_1
XFILLER_188_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _03924_ _05496_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__xnor2_1
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18256_ _01954_ _01955_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__nand2_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15468_ _08084_ _08112_ _08103_ vssd1 vssd1 vccd1 vccd1 _08113_ sky130_fd_sc_hd__or3_1
XFILLER_129_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17207_ _09783_ _09787_ _09788_ vssd1 vssd1 vccd1 vccd1 _09790_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14419_ _07154_ _07155_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__or2_1
X_18187_ _01885_ _01886_ _01876_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__a21o_1
XFILLER_156_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15399_ rbzero.wall_tracer.visualWallDist\[1\] _07925_ vssd1 vssd1 vccd1 vccd1 _08044_
+ sky130_fd_sc_hd__nand2_4
XFILLER_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17138_ _07524_ _09763_ rbzero.row_render.size\[1\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00529_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17069_ _09707_ _09708_ vssd1 vssd1 vccd1 vccd1 _09709_ sky130_fd_sc_hd__xnor2_4
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20982_ clknet_leaf_11_i_clk _00751_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21603_ net144 _01372_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[54\] sky130_fd_sc_hd__dfxtp_1
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21534_ net455 _01303_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21465_ net386 _01234_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20416_ _03272_ _03325_ _03326_ _03327_ rbzero.texV\[-12\] vssd1 vssd1 vccd1 vccd1
+ _01384_ sky130_fd_sc_hd__a32o_1
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21396_ net317 _01165_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11080_ _03890_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ _07503_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11982_ rbzero.tex_b1\[13\] rbzero.tex_b1\[12\] _04291_ vssd1 vssd1 vccd1 vccd1 _04757_
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13721_ _06427_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__or2b_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10933_ _03813_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_72_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16440_ _07970_ vssd1 vssd1 vccd1 vccd1 _09085_ sky130_fd_sc_hd__buf_4
X_10864_ _03777_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__clkbuf_1
X_13652_ _05824_ _06080_ _06282_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__o21ai_1
XFILLER_72_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12603_ rbzero.debug_overlay.facingY\[-6\] rbzero.wall_tracer.rayAddendY\[2\] vssd1
+ vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__nand2_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _09013_ _09015_ vssd1 vssd1 vccd1 vccd1 _09016_ sky130_fd_sc_hd__nor2_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _03741_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__clkbuf_1
X_13583_ _06316_ _06318_ _06319_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__a21o_1
XFILLER_24_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18110_ _01807_ _01810_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__nand2_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _07966_ vssd1 vssd1 vccd1 vccd1 _07967_ sky130_fd_sc_hd__clkbuf_4
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _02678_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__clkbuf_1
X_12534_ rbzero.debug_overlay.facingY\[-1\] rbzero.wall_tracer.rayAddendY\[7\] _05286_
+ _05287_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__a31o_1
XFILLER_157_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18041_ _01741_ _01742_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__xnor2_2
X_15253_ rbzero.debug_overlay.playerX\[-6\] _07897_ vssd1 vssd1 vccd1 vccd1 _07898_
+ sky130_fd_sc_hd__or2_2
XFILLER_184_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12465_ rbzero.wall_tracer.trackDistY\[6\] vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__inv_2
Xtop_ew_algofoogle_90 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_90/HI zeros[0] sky130_fd_sc_hd__conb_1
XFILLER_172_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14204_ _06704_ _06690_ _06663_ _05825_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__o22a_1
XFILLER_158_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11416_ gpout0.hpos\[3\] _04189_ _04187_ _04022_ _04195_ vssd1 vssd1 vccd1 vccd1
+ _04196_ sky130_fd_sc_hd__a221o_1
X_12396_ net68 _05142_ _05161_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__a211o_1
X_15184_ _07800_ _07812_ _07814_ vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__a21o_1
XFILLER_153_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ _06861_ _06871_ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__nor2_1
XFILLER_99_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11347_ _04084_ _04087_ _04114_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a21oi_1
X_19992_ rbzero.pov.ready_buffer\[18\] _03246_ _03248_ rbzero.debug_overlay.vplaneX\[-2\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__a221o_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14066_ _06787_ _06791_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__xnor2_1
X_18943_ rbzero.pov.spi_buffer\[5\] rbzero.pov.ready_buffer\[5\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02601_ sky130_fd_sc_hd__mux2_1
XFILLER_98_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11278_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] vssd1 vssd1
+ vccd1 vccd1 _04058_ sky130_fd_sc_hd__or2_1
XFILLER_141_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13017_ _05700_ _05731_ _05746_ _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__and4bb_2
X_18874_ _02537_ _02539_ _02538_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a21boi_1
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17825_ _10126_ _01528_ _10271_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__a21oi_1
XFILLER_121_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1 rbzero.tex_r1\[40\] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17756_ _09368_ _09703_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__nand2_1
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14968_ rbzero.wall_tracer.stepDistX\[-9\] _07502_ _07650_ vssd1 vssd1 vccd1 vccd1
+ _07654_ sky130_fd_sc_hd__mux2_1
XFILLER_207_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16707_ _09265_ _09240_ vssd1 vssd1 vccd1 vccd1 _09349_ sky130_fd_sc_hd__or2b_1
X_13919_ _06639_ _06654_ _06655_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17687_ _10243_ _10251_ vssd1 vssd1 vccd1 vccd1 _10252_ sky130_fd_sc_hd__xnor2_2
X_14899_ _07591_ _07606_ _07607_ _04039_ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__o211a_1
X_19426_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.debug_overlay.vplaneY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__and2_1
X_16638_ _09278_ _09280_ vssd1 vssd1 vccd1 vccd1 _09281_ sky130_fd_sc_hd__xor2_1
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19357_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__or2_1
XFILLER_204_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16569_ _08160_ _09165_ _09211_ vssd1 vssd1 vccd1 vccd1 _09212_ sky130_fd_sc_hd__or3b_1
XFILLER_200_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18308_ _01817_ _01896_ _02007_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a21oi_1
XFILLER_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19288_ _02792_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__inv_2
XFILLER_198_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18239_ _10239_ _09027_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__nor2_2
XFILLER_198_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21250_ clknet_leaf_86_i_clk _01019_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_8_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21181_ clknet_leaf_7_i_clk _00950_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20965_ clknet_leaf_5_i_clk _00734_ vssd1 vssd1 vccd1 vccd1 rbzero.othery\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ clknet_leaf_85_i_clk _00665_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10580_ rbzero.tex_r0\[1\] rbzero.tex_r0\[0\] _03624_ vssd1 vssd1 vccd1 vccd1 _03628_
+ sky130_fd_sc_hd__mux2_1
XFILLER_142_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21517_ net438 _01286_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_167_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12250_ _04984_ _04995_ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__or3b_2
XFILLER_182_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21448_ net369 _01217_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11201_ rbzero.map_rom.f1 _03942_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__nand2_1
XFILLER_108_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12181_ _04907_ _04949_ _04951_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__a21oi_1
XFILLER_163_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21379_ net300 _01148_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11132_ rbzero.map_rom.a6 vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__inv_2
XFILLER_134_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19627__79 clknet_1_0__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__inv_2
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15940_ _08539_ _08541_ vssd1 vssd1 vccd1 vccd1 _08585_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11063_ _03881_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15871_ _08199_ _08201_ _08515_ vssd1 vssd1 vccd1 vccd1 _08516_ sky130_fd_sc_hd__and3_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17610_ _10174_ _10175_ _10031_ _10033_ vssd1 vssd1 vccd1 vccd1 _10176_ sky130_fd_sc_hd__a211o_1
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14822_ _07486_ _07455_ _07548_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__a21oi_4
XFILLER_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ _02252_ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__xor2_1
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _10098_ _10106_ vssd1 vssd1 vccd1 vccd1 _10107_ sky130_fd_sc_hd__xnor2_2
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _07486_ vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__buf_4
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ rbzero.tex_b1\[17\] rbzero.tex_b1\[16\] _04356_ vssd1 vssd1 vccd1 vccd1 _04740_
+ sky130_fd_sc_hd__mux2_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _06405_ _06410_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__xor2_1
XFILLER_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17472_ _09614_ _10022_ vssd1 vssd1 vccd1 vccd1 _10038_ sky130_fd_sc_hd__nand2_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10916_ _03804_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__clkbuf_1
X_14684_ _07419_ _07420_ _05741_ _07106_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__a211o_1
XFILLER_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11896_ rbzero.tex_b0\[11\] _04327_ _04328_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__and3_1
XFILLER_204_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19211_ rbzero.spi_registers.new_floor\[1\] rbzero.spi_registers.got_new_floor _02711_
+ _03911_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__a31o_1
X_16423_ _09067_ _08955_ vssd1 vssd1 vccd1 vccd1 _09068_ sky130_fd_sc_hd__xnor2_4
X_13635_ _06350_ _06370_ _06371_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__o21a_1
X_10847_ _03768_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_160_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19142_ rbzero.spi_registers.got_new_other _02708_ vssd1 vssd1 vccd1 vccd1 _02709_
+ sky130_fd_sc_hd__and2_1
X_16354_ _08363_ _08364_ vssd1 vssd1 vccd1 vccd1 _08999_ sky130_fd_sc_hd__nor2_1
XFILLER_13_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13566_ _06131_ _06142_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__xnor2_1
XFILLER_185_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10778_ _03732_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15305_ _07948_ _07949_ _05496_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__mux2_1
XFILLER_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19073_ rbzero.pov.spi_buffer\[67\] rbzero.pov.ready_buffer\[67\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02669_ sky130_fd_sc_hd__mux2_1
X_12517_ _05263_ rbzero.wall_tracer.trackDistY\[-4\] _05252_ rbzero.wall_tracer.trackDistX\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__a2bb2o_1
X_16285_ _08922_ _08927_ _08928_ _08929_ vssd1 vssd1 vccd1 vccd1 _08930_ sky130_fd_sc_hd__o211a_1
XFILLER_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13497_ _06209_ _06223_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__and2b_1
X_18024_ _01716_ _01724_ _01725_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__or3_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15236_ rbzero.wall_tracer.rayAddendX\[8\] rbzero.wall_tracer.rayAddendX\[7\] _05448_
+ _07821_ vssd1 vssd1 vccd1 vccd1 _07885_ sky130_fd_sc_hd__or4b_1
X_12448_ rbzero.wall_tracer.state\[1\] vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__buf_6
XFILLER_172_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ rbzero.wall_tracer.rayAddendX\[4\] rbzero.wall_tracer.rayAddendX\[3\] _07821_
+ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12379_ _05143_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__clkbuf_4
XFILLER_113_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14118_ _06848_ _06850_ _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15098_ _07742_ rbzero.wall_tracer.rayAddendX\[0\] vssd1 vssd1 vccd1 vccd1 _07757_
+ sky130_fd_sc_hd__or2_1
XFILLER_4_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19975_ rbzero.pov.ready_buffer\[26\] _03247_ _03249_ rbzero.debug_overlay.facingY\[-5\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__a221o_1
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14049_ _06742_ _06785_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__xnor2_1
X_18926_ _02589_ _02557_ _02590_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__and3b_1
XFILLER_132_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18857_ _02524_ _02526_ _02525_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__a21boi_1
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17808_ _01496_ _01511_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__xor2_2
X_18788_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.stepDistY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__nor2_1
X_17739_ _10199_ _10231_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__nand2_1
X_20400__25 clknet_1_0__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__inv_2
XFILLER_63_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20145__175 clknet_1_0__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__inv_2
X_20750_ clknet_leaf_38_i_clk _00519_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19409_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__or2_1
XFILLER_91_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20681_ clknet_leaf_45_i_clk _00465_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_189_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21302_ net223 _01071_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21233_ clknet_leaf_18_i_clk _01002_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20310__323 clknet_1_0__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__inv_2
X_21164_ clknet_leaf_89_i_clk _00933_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21095_ net185 _00864_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[35\] sky130_fd_sc_hd__dfxtp_1
X_20046_ _03283_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__clkbuf_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ rbzero.tex_g0\[11\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__and3_1
X_20948_ clknet_leaf_4_i_clk _00717_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10701_ rbzero.tex_g1\[7\] rbzero.tex_g1\[8\] _03691_ vssd1 vssd1 vccd1 vccd1 _03692_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11681_ _04004_ _04419_ _04450_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__and3_2
XFILLER_201_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20879_ clknet_leaf_97_i_clk _00648_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_13420_ _05978_ _05942_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__nor2_1
XFILLER_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10632_ _03655_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_179_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10563_ rbzero.tex_r0\[9\] rbzero.tex_r0\[8\] _03613_ vssd1 vssd1 vccd1 vccd1 _03619_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13351_ _06082_ _06087_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__xor2_1
XFILLER_195_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12302_ _03473_ _05044_ _05046_ _04317_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__a221o_1
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16070_ _08696_ _08714_ vssd1 vssd1 vccd1 vccd1 _08715_ sky130_fd_sc_hd__nand2_1
X_10494_ rbzero.tex_r0\[42\] rbzero.tex_r0\[41\] _03580_ vssd1 vssd1 vccd1 vccd1 _03583_
+ sky130_fd_sc_hd__mux2_1
X_13282_ _06010_ _06012_ _06014_ _06018_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__a22o_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15021_ rbzero.debug_overlay.vplaneX\[-8\] rbzero.wall_tracer.rayAddendX\[-8\] vssd1
+ vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__or2_1
X_12233_ _03473_ _04814_ _04317_ _04809_ _04961_ _04960_ vssd1 vssd1 vccd1 vccd1 _05003_
+ sky130_fd_sc_hd__mux4_1
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ net38 _04907_ net8 vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__and3_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11115_ _03908_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20285__300 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__inv_2
XFILLER_150_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16972_ _08162_ _09611_ vssd1 vssd1 vccd1 vccd1 _09612_ sky130_fd_sc_hd__and2_1
XFILLER_150_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12095_ net51 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__buf_6
X_19760_ _03108_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15923_ _08566_ _08567_ vssd1 vssd1 vccd1 vccd1 _08568_ sky130_fd_sc_hd__nand2_1
X_18711_ _05532_ _02403_ _02404_ _02399_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__o31a_1
X_11046_ _03872_ vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__clkbuf_1
X_19691_ _03072_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18642_ _01620_ _09292_ _02239_ _02337_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__o31a_1
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03291_ _03291_ vssd1 vssd1 vccd1 vccd1 clknet_0__03291_ sky130_fd_sc_hd__clkbuf_16
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _08084_ _08041_ _08498_ vssd1 vssd1 vccd1 vccd1 _08499_ sky130_fd_sc_hd__or3_1
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _07511_ _07534_ vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__nor2_1
XFILLER_206_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ _02192_ _02185_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__or2b_1
XFILLER_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15785_ _08330_ _08415_ _08429_ vssd1 vssd1 vccd1 vccd1 _08430_ sky130_fd_sc_hd__and3_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12997_ _05589_ _05704_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__xor2_2
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17524_ _09963_ _09969_ _10089_ vssd1 vssd1 vccd1 vccd1 _10090_ sky130_fd_sc_hd__a21o_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14736_ _07469_ _07470_ _05952_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__mux2_1
XFILLER_189_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11948_ _04254_ _04719_ _04723_ _04371_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a211o_1
XFILLER_189_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17455_ _10019_ _10021_ vssd1 vssd1 vccd1 vccd1 _10022_ sky130_fd_sc_hd__xor2_4
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14667_ _07375_ _07403_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__nand2_1
XFILLER_177_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11879_ rbzero.tex_g1\[29\] rbzero.tex_g1\[28\] _04336_ vssd1 vssd1 vccd1 vccd1 _04656_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16406_ _08371_ _08411_ vssd1 vssd1 vccd1 vccd1 _09051_ sky130_fd_sc_hd__nor2_1
XFILLER_20_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13618_ _06311_ _06314_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__xnor2_1
X_17386_ _09920_ _09921_ _09951_ vssd1 vssd1 vccd1 vccd1 _09953_ sky130_fd_sc_hd__nand3_1
XFILLER_186_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ _07218_ _07323_ _07334_ _07332_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__a31o_1
X_19125_ _02697_ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16337_ _08218_ _08232_ _08208_ _08981_ vssd1 vssd1 vccd1 vccd1 _08982_ sky130_fd_sc_hd__a31o_1
XFILLER_119_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13549_ _05975_ _06285_ _05921_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__and3b_1
XFILLER_186_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19056_ _02593_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__buf_4
X_16268_ _08215_ _08335_ _08856_ vssd1 vssd1 vccd1 vccd1 _08913_ sky130_fd_sc_hd__a21o_1
X_18007_ _01462_ _09359_ _01707_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__o21ai_1
XFILLER_161_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15219_ _07820_ rbzero.wall_tracer.rayAddendX\[9\] vssd1 vssd1 vccd1 vccd1 _07870_
+ sky130_fd_sc_hd__nand2_1
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16199_ _08836_ _08842_ _08843_ vssd1 vssd1 vccd1 vccd1 _08844_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_i_clk clknet_opt_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19958_ _03245_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__clkbuf_4
XFILLER_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18909_ rbzero.spi_registers.spi_counter\[1\] _02576_ vssd1 vssd1 vccd1 vccd1 _02578_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_206_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19889_ _03194_ _03193_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__nand2_1
XFILLER_171_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20802_ clknet_leaf_25_i_clk _00571_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20733_ clknet_3_5_0_i_clk _00502_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20664_ clknet_leaf_63_i_clk _00448_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20595_ _02833_ _03460_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21216_ clknet_leaf_20_i_clk _00985_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_105_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21147_ clknet_leaf_88_i_clk _00916_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21078_ net168 _00847_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20029_ _09749_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__buf_4
XFILLER_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12920_ _05567_ _05575_ _05576_ _05656_ _05563_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__o2111a_1
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ rbzero.wall_tracer.visualWallDist\[-10\] rbzero.wall_tracer.rayAddendY\[-2\]
+ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__mux2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _04253_ _04575_ _04579_ _04119_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__a211o_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ rbzero.wall_tracer.visualWallDist\[-10\] _04012_ vssd1 vssd1 vccd1 vccd1
+ _08215_ sky130_fd_sc_hd__nand2_8
X_20280__296 clknet_1_1__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__inv_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12782_ rbzero.wall_tracer.mapX\[5\] _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__xnor2_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14521_ _07254_ _07257_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__xnor2_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ rbzero.debug_overlay.playerX\[5\] _04444_ _04439_ _04452_ rbzero.debug_overlay.playerX\[3\]
+ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__a32o_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17240_ _08940_ _08943_ _05204_ vssd1 vssd1 vccd1 vccd1 _09818_ sky130_fd_sc_hd__a21oi_1
XFILLER_14_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14452_ _07175_ _07180_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__xor2_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _04441_ _04442_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__nor2_1
XFILLER_202_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ _06069_ _06074_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__xor2_1
X_10615_ _03481_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__buf_4
XFILLER_31_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17171_ rbzero.traced_texa\[0\] _09768_ _09769_ rbzero.wall_tracer.visualWallDist\[0\]
+ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__a22o_1
X_14383_ _07115_ _07119_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__xnor2_1
X_20317__329 clknet_1_0__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__inv_2
X_11595_ _04140_ _04355_ _04373_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__or3_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16122_ _08284_ vssd1 vssd1 vccd1 vccd1 _08767_ sky130_fd_sc_hd__buf_4
XFILLER_31_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13334_ _06053_ _06056_ _06061_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__a21o_1
XFILLER_182_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10546_ rbzero.tex_r0\[17\] rbzero.tex_r0\[16\] _03602_ vssd1 vssd1 vccd1 vccd1 _03610_
+ sky130_fd_sc_hd__mux2_1
XFILLER_116_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16053_ _08640_ _08648_ vssd1 vssd1 vccd1 vccd1 _08698_ sky130_fd_sc_hd__xnor2_1
X_13265_ _05945_ _05949_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nand2_4
X_10477_ rbzero.tex_r0\[50\] rbzero.tex_r0\[49\] _03569_ vssd1 vssd1 vccd1 vccd1 _03574_
+ sky130_fd_sc_hd__mux2_1
XFILLER_157_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15004_ _07672_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__clkbuf_1
X_12216_ net18 _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nand2_1
XFILLER_124_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13196_ _05591_ _05740_ _05931_ _05893_ _05932_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__a41o_1
XFILLER_151_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19812_ rbzero.pov.sclk_buffer\[2\] rbzero.pov.sclk_buffer\[1\] _05189_ vssd1 vssd1
+ vccd1 vccd1 _03135_ sky130_fd_sc_hd__mux2_1
XFILLER_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12147_ _04907_ net8 vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__nor2_4
XFILLER_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03312_ clknet_0__03312_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03312_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19743_ _03099_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12078_ net4 vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__inv_2
X_16955_ _09207_ _09330_ _09457_ _09595_ vssd1 vssd1 vccd1 vccd1 _09596_ sky130_fd_sc_hd__a31o_2
XFILLER_42_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15906_ _08483_ _08480_ vssd1 vssd1 vccd1 vccd1 _08551_ sky130_fd_sc_hd__nand2_1
X_11029_ _03863_ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__clkbuf_1
X_16886_ _09526_ _08356_ _09524_ vssd1 vssd1 vccd1 vccd1 _09527_ sky130_fd_sc_hd__o21ai_1
X_19674_ _03063_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18625_ _09889_ _02321_ _09780_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__a21oi_1
X_15837_ _07912_ _08019_ _08020_ vssd1 vssd1 vccd1 vccd1 _08482_ sky130_fd_sc_hd__or3_1
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18556_ _02159_ _02143_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__or2b_1
X_15768_ _08154_ _08167_ vssd1 vssd1 vccd1 vccd1 _08413_ sky130_fd_sc_hd__or2b_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17507_ _09522_ _08159_ _08151_ _09661_ vssd1 vssd1 vccd1 vccd1 _10073_ sky130_fd_sc_hd__o22ai_1
X_14719_ _07455_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__buf_4
X_18487_ _02088_ _02090_ _02087_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a21bo_1
XFILLER_178_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15699_ _08340_ _08341_ _08342_ vssd1 vssd1 vccd1 vccd1 _08344_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17438_ _09702_ _09713_ _10004_ vssd1 vssd1 vccd1 vccd1 _10005_ sky130_fd_sc_hd__a21o_1
XFILLER_166_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 _08039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_26 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_37 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_48 _08096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ _09926_ _09935_ vssd1 vssd1 vccd1 vccd1 _09936_ sky130_fd_sc_hd__nand2_1
XANTENNA_59 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20257__276 clknet_1_0__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__inv_2
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19108_ _02687_ vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__clkbuf_1
XFILLER_146_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039_ _02651_ vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21001_ clknet_leaf_11_i_clk _00770_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20716_ clknet_leaf_72_i_clk _00006_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20647_ clknet_leaf_62_i_clk _00431_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10400_ _03531_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11380_ rbzero.row_render.size\[5\] vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__inv_2
XFILLER_176_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20578_ _03450_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_109_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10331_ _03495_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13050_ _05695_ _05702_ _05785_ _05786_ _05766_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__o311a_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12001_ rbzero.tex_b1\[53\] rbzero.tex_b1\[52\] _04212_ vssd1 vssd1 vccd1 vccd1 _04776_
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16740_ _09348_ _09381_ vssd1 vssd1 vccd1 vccd1 _09382_ sky130_fd_sc_hd__xnor2_1
X_13952_ _06245_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__clkbuf_4
XFILLER_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12903_ _05615_ _05639_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__xor2_2
XFILLER_98_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16671_ _09113_ _09152_ _09313_ vssd1 vssd1 vccd1 vccd1 _09314_ sky130_fd_sc_hd__a21o_1
X_13883_ _06239_ _06245_ _06202_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__or3_1
XFILLER_189_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18410_ _01946_ _01949_ _02108_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a21oi_4
X_15622_ _07981_ _08177_ _08266_ _08264_ vssd1 vssd1 vccd1 vccd1 _08267_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19390_ rbzero.wall_tracer.rayAddendY\[-1\] _07706_ _02876_ _07703_ vssd1 vssd1 vccd1
+ vccd1 _02877_ sky130_fd_sc_hd__a22o_1
X_12834_ _05570_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__buf_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _10238_ _09294_ _09977_ _01737_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__o22ai_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _08171_ _08197_ _05193_ vssd1 vssd1 vccd1 vccd1 _08198_ sky130_fd_sc_hd__o21ai_1
XFILLER_188_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _03936_ _05503_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__nor2_1
XFILLER_199_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14504_ _06239_ _07071_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__nor2_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18272_ _01968_ _01971_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__xnor2_1
X_11716_ rbzero.debug_overlay.facingX\[-5\] _04454_ _04455_ rbzero.debug_overlay.facingX\[-7\]
+ _04494_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__a221o_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15484_ _08035_ vssd1 vssd1 vccd1 vccd1 _08129_ sky130_fd_sc_hd__clkbuf_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12696_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__nor2_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17223_ rbzero.wall_tracer.mapX\[11\] _09781_ _09779_ _09802_ vssd1 vssd1 vccd1 vccd1
+ _00576_ sky130_fd_sc_hd__a22o_1
XFILLER_147_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14435_ _07171_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__dlymetal6s2s_1
X_11647_ _04005_ _04023_ _04425_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__a21o_2
XFILLER_128_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 i_gpout1_sel[5] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_6
XFILLER_174_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17154_ rbzero.row_render.texu\[4\] _09766_ _07728_ rbzero.wall_tracer.texu\[4\]
+ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__a22o_1
Xinput24 i_gpout3_sel[4] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_6
XFILLER_196_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput35 i_gpout5_sel[3] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_4
XFILLER_155_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14366_ _05793_ _07041_ _07102_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__a21oi_1
Xinput46 i_tex_in[0] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__buf_4
X_11578_ rbzero.tex_r1\[19\] rbzero.tex_r1\[18\] _04356_ vssd1 vssd1 vccd1 vccd1 _04357_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16105_ _08744_ _08749_ vssd1 vssd1 vccd1 vccd1 _08750_ sky130_fd_sc_hd__xor2_1
XFILLER_116_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13317_ _05939_ _05961_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__nor2_1
X_10529_ rbzero.tex_r0\[25\] rbzero.tex_r0\[24\] _03591_ vssd1 vssd1 vccd1 vccd1 _03601_
+ sky130_fd_sc_hd__mux2_1
X_17085_ _09722_ _09724_ vssd1 vssd1 vccd1 vccd1 _09725_ sky130_fd_sc_hd__xor2_2
XFILLER_7_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14297_ _07031_ _07033_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__xor2_2
XFILLER_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16036_ _08624_ _08628_ vssd1 vssd1 vccd1 vccd1 _08681_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13248_ _05983_ _05975_ _05984_ _05974_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__o22a_1
XFILLER_170_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _05695_ _05677_ _05801_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__mux2_1
XFILLER_97_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_17987_ _09249_ _01576_ _01579_ _01577_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__o22a_1
XFILLER_42_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19726_ _03090_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__clkbuf_1
X_16938_ _09538_ _09578_ vssd1 vssd1 vccd1 vccd1 _09579_ sky130_fd_sc_hd__xnor2_1
XFILLER_42_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19657_ _03054_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16869_ _09507_ _09509_ vssd1 vssd1 vccd1 vccd1 _09510_ sky130_fd_sc_hd__nor2_1
XFILLER_77_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19596__51 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__inv_2
X_18608_ _02303_ _02304_ vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_95_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18539_ _02149_ _02156_ _02155_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__o21bai_1
XFILLER_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21550_ net471 _01319_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20501_ _03398_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__inv_2
X_21481_ net402 _01250_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20432_ _03333_ _03334_ _03335_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__o21ai_1
XFILLER_107_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20294_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__buf_1
XFILLER_134_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10880_ rbzero.tex_b1\[50\] rbzero.tex_b1\[51\] _03784_ vssd1 vssd1 vccd1 vccd1 _03786_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12550_ rbzero.debug_overlay.facingY\[-4\] rbzero.wall_tracer.rayAddendY\[4\] vssd1
+ vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__nor2_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11501_ _04230_ _04276_ _04280_ _04232_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__a211o_1
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ rbzero.wall_tracer.trackDistX\[-5\] vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__inv_2
XFILLER_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03315_ clknet_0__03315_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03315_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_156_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14220_ _06923_ _06931_ _06956_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__a21boi_1
X_11432_ _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__buf_4
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _05825_ _06678_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__nor2_1
X_11363_ _04100_ _04114_ _04120_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__nor3_4
XFILLER_192_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13102_ _05710_ _05713_ _05715_ _05687_ _05791_ _05826_ vssd1 vssd1 vccd1 vccd1 _05839_
+ sky130_fd_sc_hd__mux4_1
X_10314_ _03486_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__clkbuf_1
X_14082_ _06685_ _06695_ _06702_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__and3_1
XFILLER_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11294_ rbzero.texV\[4\] _04072_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__a21boi_1
XFILLER_4_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17910_ _01502_ _01510_ _01612_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__a21o_1
X_13033_ _05719_ _05721_ _05734_ _05708_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__or4_1
XFILLER_156_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18890_ rbzero.spi_registers.spi_cmd\[3\] rbzero.spi_registers.spi_cmd\[2\] vssd1
+ vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__nor2_1
XFILLER_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17841_ _10195_ _10284_ _01544_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__a21oi_1
XFILLER_120_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17772_ _08149_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__clkbuf_4
XFILLER_19_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14984_ _00008_ _07549_ _07662_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__a21oi_1
X_19511_ _02905_ rbzero.wall_tracer.rayAddendY\[8\] vssd1 vssd1 vccd1 vccd1 _02989_
+ sky130_fd_sc_hd__xnor2_1
X_16723_ _09243_ _08821_ _08419_ vssd1 vssd1 vccd1 vccd1 _09365_ sky130_fd_sc_hd__or3_1
X_13935_ _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__clkbuf_4
XFILLER_93_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16654_ _09291_ _09293_ _09296_ vssd1 vssd1 vccd1 vccd1 _09297_ sky130_fd_sc_hd__nand3_1
XFILLER_19_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19442_ _02921_ _02922_ _02923_ _02924_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__a211oi_2
X_13866_ _06602_ _06557_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__xor2_4
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03042_ _03042_ vssd1 vssd1 vccd1 vccd1 clknet_0__03042_ sky130_fd_sc_hd__clkbuf_16
X_15605_ _07945_ _08238_ vssd1 vssd1 vccd1 vccd1 _08250_ sky130_fd_sc_hd__nor2_4
XFILLER_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12817_ _05548_ _05552_ _05554_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__or3_1
X_16585_ _08329_ _08427_ vssd1 vssd1 vccd1 vccd1 _09228_ sky130_fd_sc_hd__nor2_1
XFILLER_50_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19373_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.wall_tracer.rayAddendY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__nand2_1
XFILLER_90_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13797_ _06529_ _06533_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__nand2_1
XFILLER_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18324_ _01902_ _02012_ _02011_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__a21o_1
X_15536_ _07560_ _07562_ _08171_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__or3_1
XFILLER_163_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__buf_4
XFILLER_203_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18255_ _08257_ _01475_ _01476_ _01739_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__o22ai_1
X_15467_ _08102_ vssd1 vssd1 vccd1 vccd1 _08112_ sky130_fd_sc_hd__clkbuf_4
XFILLER_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12679_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__nand2_1
XFILLER_175_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17206_ _09783_ _09787_ _09788_ vssd1 vssd1 vccd1 vccd1 _09789_ sky130_fd_sc_hd__or3_1
XFILLER_200_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14418_ _07146_ _07153_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__nor2_1
X_18186_ _01876_ _01885_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__nand3_1
XFILLER_191_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15398_ _08035_ _08042_ vssd1 vssd1 vccd1 vccd1 _08043_ sky130_fd_sc_hd__or2_1
XFILLER_144_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17137_ _07514_ _09763_ rbzero.row_render.size\[0\] _09764_ vssd1 vssd1 vccd1 vccd1
+ _00528_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_155_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14349_ _07084_ _07085_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__nand2_1
XFILLER_156_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17068_ _08519_ _09565_ vssd1 vssd1 vccd1 vccd1 _09708_ sky130_fd_sc_hd__or2_2
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16019_ _08622_ _08653_ vssd1 vssd1 vccd1 vccd1 _08664_ sky130_fd_sc_hd__nor2_1
XFILLER_135_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20369__377 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__inv_2
XFILLER_97_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20068__105 clknet_1_0__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__inv_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19709_ rbzero.pov.spi_buffer\[29\] rbzero.pov.spi_buffer\[30\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03082_ sky130_fd_sc_hd__mux2_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20981_ clknet_leaf_11_i_clk _00750_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03309_ _03309_ vssd1 vssd1 vccd1 vccd1 clknet_0__03309_ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21602_ net143 _01371_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[53\] sky130_fd_sc_hd__dfxtp_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_13_0_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_13_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21533_ net454 _01302_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21464_ net385 _01233_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20415_ _02695_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__buf_4
XFILLER_193_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21395_ net316 _01164_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ rbzero.tex_b1\[15\] _04221_ _04222_ _04218_ vssd1 vssd1 vccd1 vccd1 _04756_
+ sky130_fd_sc_hd__a31o_1
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13720_ _06438_ _06455_ _06456_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10932_ rbzero.tex_b1\[25\] rbzero.tex_b1\[26\] _03806_ vssd1 vssd1 vccd1 vccd1 _03813_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19575__32 clknet_1_1__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__inv_2
XFILLER_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13651_ _05988_ _06380_ _06387_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__o21bai_1
XFILLER_44_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10863_ rbzero.tex_b1\[58\] rbzero.tex_b1\[59\] _03773_ vssd1 vssd1 vccd1 vccd1 _03777_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12602_ rbzero.wall_tracer.rayAddendY\[-4\] rbzero.wall_tracer.rayAddendY\[-3\] rbzero.wall_tracer.rayAddendY\[-2\]
+ _05355_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__or4_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _08361_ _07967_ _08097_ _09014_ vssd1 vssd1 vccd1 vccd1 _09015_ sky130_fd_sc_hd__o31a_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13582_ _06309_ _06315_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__nor2_1
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ rbzero.tex_g0\[28\] rbzero.tex_g0\[27\] _03740_ vssd1 vssd1 vccd1 vccd1 _03741_
+ sky130_fd_sc_hd__mux2_1
XFILLER_197_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19590__46 clknet_1_0__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__inv_2
XFILLER_185_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _07964_ _07965_ vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__or2_1
XFILLER_9_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__and2_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18040_ _08257_ _01620_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__nor2_1
X_15252_ rbzero.debug_overlay.playerX\[-7\] rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__or3_1
X_12464_ _05217_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.trackDistY\[7\]
+ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__a22o_1
XFILLER_200_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_80 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_80/HI o_rgb[10] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_91 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_91/HI zeros[1] sky130_fd_sc_hd__conb_1
XFILLER_184_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14203_ _05825_ _06690_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__nor2_1
X_11415_ gpout0.hpos\[3\] _04189_ _04191_ _04194_ vssd1 vssd1 vccd1 vccd1 _04195_
+ sky130_fd_sc_hd__o211a_1
X_15183_ _07835_ _07836_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__nand2_1
X_12395_ net47 _05145_ _05143_ _05149_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__a31o_1
XFILLER_158_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14134_ _06862_ _06869_ _06870_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__a21boi_1
XFILLER_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11346_ _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__buf_4
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19991_ rbzero.pov.ready_buffer\[17\] _03252_ _03253_ _04462_ _03254_ vssd1 vssd1
+ vccd1 vccd1 _01032_ sky130_fd_sc_hd__o221a_1
XFILLER_67_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14065_ _06713_ _06801_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__and2_1
X_18942_ _02600_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__clkbuf_1
X_11277_ rbzero.traced_texVinit\[7\] rbzero.spi_registers.vshift\[4\] vssd1 vssd1
+ vccd1 vccd1 _04057_ sky130_fd_sc_hd__nand2_1
XFILLER_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13016_ _05747_ _05684_ _05749_ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__o211a_1
X_18873_ _02544_ _02545_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__nand2_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17824_ _01526_ _01527_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__xor2_1
XFILLER_0_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2 rbzero.pov.ready_buffer\[31\] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_181_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17755_ _09249_ _10200_ _01458_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__o21ba_1
XFILLER_130_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14967_ _07653_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16706_ _09222_ _09236_ _09234_ vssd1 vssd1 vccd1 vccd1 _09348_ sky130_fd_sc_hd__a21o_1
X_12063__1 clknet_1_1__leaf__04835_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__inv_2
X_13918_ _06617_ _06638_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__and2_1
X_17686_ _10247_ _10250_ vssd1 vssd1 vccd1 vccd1 _10251_ sky130_fd_sc_hd__xor2_2
X_14898_ rbzero.wall_tracer.visualWallDist\[-8\] _07595_ vssd1 vssd1 vccd1 vccd1 _07607_
+ sky130_fd_sc_hd__or2_1
XFILLER_39_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19425_ _02893_ _02896_ _02907_ _07676_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a31o_1
XFILLER_90_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16637_ _08237_ _09279_ _08170_ vssd1 vssd1 vccd1 vccd1 _09280_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13849_ _06574_ _06585_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__nand2_1
XFILLER_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19356_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__nand2_1
X_16568_ _08054_ _09029_ vssd1 vssd1 vccd1 vccd1 _09211_ sky130_fd_sc_hd__nor2_1
XFILLER_204_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18307_ _01892_ _01893_ _01895_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__and3_1
XFILLER_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15519_ _08161_ _08163_ vssd1 vssd1 vccd1 vccd1 _08164_ sky130_fd_sc_hd__nor2_1
X_16499_ _08979_ _08239_ _09141_ _09142_ vssd1 vssd1 vccd1 vccd1 _09143_ sky130_fd_sc_hd__o31a_1
X_19287_ _02798_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18238_ _01936_ _01937_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__xor2_2
XFILLER_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18169_ _01868_ _01869_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__xnor2_1
XFILLER_156_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21180_ clknet_leaf_7_i_clk _00949_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20964_ clknet_leaf_5_i_clk _00733_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20895_ clknet_leaf_68_i_clk _00664_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20122__154 clknet_1_1__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__inv_2
XFILLER_142_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21516_ net437 _01285_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_127_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21447_ net368 _01216_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11200_ _03936_ _03982_ rbzero.map_rom.a6 rbzero.map_rom.f2 vssd1 vssd1 vccd1 vccd1
+ _03989_ sky130_fd_sc_hd__a22o_1
X_12180_ net9 _04950_ net11 vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__a21bo_1
XFILLER_181_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21378_ net299 _01147_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11131_ rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__inv_2
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11062_ rbzero.tex_b0\[28\] rbzero.tex_b0\[27\] _03876_ vssd1 vssd1 vccd1 vccd1 _03881_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15870_ rbzero.wall_tracer.visualWallDist\[-12\] _07925_ vssd1 vssd1 vccd1 vccd1
+ _08515_ sky130_fd_sc_hd__and2_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14821_ _05834_ _07392_ _07472_ _07527_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__a22o_1
XFILLER_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17540_ _10103_ _10105_ vssd1 vssd1 vccd1 vccd1 _10106_ sky130_fd_sc_hd__xor2_2
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _05834_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__buf_4
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ rbzero.tex_b1\[19\] rbzero.tex_b1\[18\] _04356_ vssd1 vssd1 vccd1 vccd1 _04739_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _06431_ _06433_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__xor2_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ _10019_ _10021_ vssd1 vssd1 vccd1 vccd1 _10037_ sky130_fd_sc_hd__or2_1
X_10915_ rbzero.tex_b1\[33\] rbzero.tex_b1\[34\] _03795_ vssd1 vssd1 vccd1 vccd1 _03804_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14683_ _07107_ _07413_ _07414_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__or3_2
X_11895_ rbzero.tex_b0\[9\] rbzero.tex_b0\[8\] _04272_ vssd1 vssd1 vccd1 vccd1 _04671_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19210_ _02753_ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__clkbuf_1
X_13634_ _06351_ _06369_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__nand2_1
XFILLER_60_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16422_ _08617_ _08672_ vssd1 vssd1 vccd1 vccd1 _09067_ sky130_fd_sc_hd__xor2_2
X_10846_ rbzero.tex_g0\[3\] rbzero.tex_g0\[2\] _03762_ vssd1 vssd1 vccd1 vccd1 _03768_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16353_ _08995_ _08997_ vssd1 vssd1 vccd1 vccd1 _08998_ sky130_fd_sc_hd__xor2_4
X_19141_ _02707_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__buf_4
XFILLER_201_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13565_ _06281_ _06283_ _06301_ _06300_ _06284_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__o32a_1
X_10777_ rbzero.tex_g0\[36\] rbzero.tex_g0\[35\] _03729_ vssd1 vssd1 vccd1 vccd1 _03732_
+ sky130_fd_sc_hd__mux2_1
X_20097__131 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__inv_2
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15304_ rbzero.debug_overlay.playerX\[-4\] vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__inv_2
XFILLER_200_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19072_ _02668_ vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__clkbuf_1
X_12516_ _05261_ _05262_ _05266_ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__or4b_1
X_16284_ _08870_ _08887_ vssd1 vssd1 vccd1 vccd1 _08929_ sky130_fd_sc_hd__xnor2_1
XFILLER_146_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13496_ _06229_ _06227_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__or2b_1
XFILLER_200_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18023_ _01717_ _01619_ _01723_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__and3_1
X_15235_ rbzero.wall_tracer.rayAddendX\[10\] _07855_ _07880_ _07884_ vssd1 vssd1 vccd1
+ vccd1 _00506_ sky130_fd_sc_hd__a211o_1
X_12447_ _05202_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15166_ _07820_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__clkbuf_4
X_12378_ net33 vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__clkbuf_4
X_14117_ _06851_ _06853_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__and2b_1
X_11329_ _04048_ _04051_ _04053_ _04056_ _04108_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__a221o_1
XFILLER_10_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19974_ rbzero.pov.ready_buffer\[25\] _03247_ _03249_ rbzero.debug_overlay.facingY\[-6\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__a221o_1
X_15097_ _07678_ vssd1 vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__buf_6
XFILLER_125_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14048_ _06666_ _06708_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__nor2_1
X_18925_ rbzero.spi_registers.spi_counter\[4\] rbzero.spi_registers.spi_counter\[3\]
+ _02580_ rbzero.spi_registers.spi_counter\[5\] vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a31o_1
XFILLER_80_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18856_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.stepDistY\[8\] vssd1
+ vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__and2_1
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17807_ _01502_ _01510_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__xnor2_2
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20397__22 clknet_1_1__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__inv_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18787_ rbzero.wall_tracer.trackDistY\[-2\] _02406_ _02471_ vssd1 vssd1 vccd1 vccd1
+ _00611_ sky130_fd_sc_hd__o21ba_1
X_15999_ _08642_ _08643_ vssd1 vssd1 vccd1 vccd1 _08644_ sky130_fd_sc_hd__xnor2_2
XFILLER_94_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17738_ _10042_ _10194_ _10192_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__a21o_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17669_ _10103_ _10105_ vssd1 vssd1 vccd1 vccd1 _10234_ sky130_fd_sc_hd__nor2_1
XFILLER_51_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19408_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[1\] vssd1
+ vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__nand2_1
XFILLER_90_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20680_ clknet_leaf_44_i_clk _00464_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[9\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19339_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__nand2_1
XFILLER_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21301_ net222 _01070_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21232_ clknet_leaf_19_i_clk _01001_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_102_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21163_ clknet_leaf_87_i_clk _00932_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21094_ net184 _00863_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20045_ _03281_ _05190_ _03282_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__and3b_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ clknet_leaf_4_i_clk _00716_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _03646_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__clkbuf_4
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _04436_ _04448_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__nor2_4
X_20878_ clknet_leaf_96_i_clk _00647_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_198_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ rbzero.tex_g1\[40\] rbzero.tex_g1\[41\] _03647_ vssd1 vssd1 vccd1 vccd1 _03655_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13350_ _06083_ _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__xnor2_1
XFILLER_194_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10562_ _03618_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _04163_ _05043_ _05049_ _04809_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a22o_1
XFILLER_155_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ _06010_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__nor2_1
XFILLER_6_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10493_ _03582_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15020_ rbzero.debug_overlay.vplaneX\[-9\] rbzero.wall_tracer.rayAddendX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__nand2_1
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12232_ _04996_ _04998_ _05000_ _05001_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__o211a_2
XFILLER_182_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12163_ _04809_ _04907_ _04909_ net10 _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__o311a_1
X_11114_ rbzero.tex_b0\[3\] rbzero.tex_b0\[2\] _03898_ vssd1 vssd1 vccd1 vccd1 _03908_
+ sky130_fd_sc_hd__mux2_1
XFILLER_116_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12094_ _04851_ _04863_ _04864_ _04865_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a22o_1
X_16971_ _05211_ _09610_ vssd1 vssd1 vccd1 vccd1 _09611_ sky130_fd_sc_hd__nor2_2
XFILLER_123_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18710_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.stepDistY\[-12\]
+ _02401_ _02402_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a22oi_1
X_15922_ _08557_ _08563_ _08565_ vssd1 vssd1 vccd1 vccd1 _08567_ sky130_fd_sc_hd__nand3_1
X_11045_ rbzero.tex_b0\[36\] rbzero.tex_b0\[35\] _03865_ vssd1 vssd1 vccd1 vccd1 _03872_
+ sky130_fd_sc_hd__mux2_1
X_19690_ rbzero.pov.spi_buffer\[20\] rbzero.pov.spi_buffer\[21\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03072_ sky130_fd_sc_hd__mux2_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18641_ _02237_ _02238_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__nand2_1
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__03290_ _03290_ vssd1 vssd1 vccd1 vccd1 clknet_0__03290_ sky130_fd_sc_hd__clkbuf_16
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ _08074_ _08125_ vssd1 vssd1 vccd1 vccd1 _08498_ sky130_fd_sc_hd__or2_1
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804_ _07104_ _07450_ _05742_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__mux2_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18572_ _02039_ _02042_ _02191_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__a21o_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ _08426_ _08428_ vssd1 vssd1 vccd1 vccd1 _08429_ sky130_fd_sc_hd__nand2_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12996_ _05721_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__inv_2
XFILLER_188_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _09967_ _09968_ vssd1 vssd1 vccd1 vccd1 _10089_ sky130_fd_sc_hd__nor2_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11947_ _04225_ _04720_ _04721_ _04722_ _04208_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__o221a_1
XFILLER_18_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14735_ _07380_ _07427_ vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__nand2_1
XFILLER_73_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_999 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17454_ _09616_ _09729_ _10020_ vssd1 vssd1 vccd1 vccd1 _10021_ sky130_fd_sc_hd__a21oi_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14666_ _07400_ _07402_ _05892_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__mux2_1
XFILLER_177_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11878_ _04653_ _04654_ _04265_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__mux2_1
XFILLER_162_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16405_ _09025_ _09049_ vssd1 vssd1 vccd1 vccd1 _09050_ sky130_fd_sc_hd__xnor2_4
X_13617_ _06353_ _06318_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__xnor2_1
XFILLER_189_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10829_ rbzero.tex_g0\[11\] rbzero.tex_g0\[10\] _03751_ vssd1 vssd1 vccd1 vccd1 _03759_
+ sky130_fd_sc_hd__mux2_1
X_17385_ _09920_ _09921_ _09951_ vssd1 vssd1 vccd1 vccd1 _09952_ sky130_fd_sc_hd__a21o_1
XFILLER_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14597_ _07332_ _07333_ vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__nor2_1
X_19124_ rbzero.spi_registers.mosi rbzero.spi_registers.mosi_buffer\[0\] _05189_ vssd1
+ vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__mux2_1
XFILLER_201_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16336_ _07571_ vssd1 vssd1 vccd1 vccd1 _08981_ sky130_fd_sc_hd__inv_2
X_13548_ _05945_ _05949_ _05990_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__a21oi_1
XFILLER_201_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16267_ _08226_ _08816_ _08162_ _08160_ vssd1 vssd1 vccd1 vccd1 _08912_ sky130_fd_sc_hd__or4_1
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19055_ _02659_ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_145_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13479_ _05990_ _06080_ _06084_ _05991_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__o22a_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18006_ _09522_ _09217_ _01707_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__or3_1
X_15218_ rbzero.wall_tracer.rayAddendX\[8\] rbzero.wall_tracer.rayAddendX\[7\] _07821_
+ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__o21a_1
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16198_ _08815_ _08835_ vssd1 vssd1 vccd1 vccd1 _08843_ sky130_fd_sc_hd__nor2_1
XFILLER_126_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _07791_ _07793_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__and2_1
XFILLER_142_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19957_ rbzero.pov.ready _02707_ _02820_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__and3_1
X_20151__180 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__inv_2
XFILLER_68_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18908_ _02577_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19888_ _03194_ rbzero.pov.ready_buffer\[44\] _02822_ vssd1 vssd1 vccd1 vccd1 _03195_
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18839_ _02516_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20801_ clknet_leaf_44_i_clk _00570_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20732_ clknet_leaf_68_i_clk _00501_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20663_ clknet_leaf_62_i_clk _00447_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20594_ _02828_ _02834_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__and2b_1
XFILLER_177_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_4_0_i_clk clknet_2_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_136_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20234__255 clknet_1_0__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__inv_2
XFILLER_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21215_ clknet_leaf_20_i_clk _00984_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_133_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21146_ clknet_leaf_88_i_clk _00915_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21077_ net167 _00846_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20028_ _02704_ _03270_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__nor2_1
XFILLER_150_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ _04000_ _05472_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__and2_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _04224_ _04576_ _04577_ _04578_ _04141_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__o221a_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _05512_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__clkbuf_4
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ _07256_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__inv_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ rbzero.debug_overlay.playerX\[1\] _04449_ _04464_ rbzero.debug_overlay.playerX\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__a22o_1
X_20391__17 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__inv_2
XFILLER_148_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14451_ _06704_ _06761_ _07060_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__o21ba_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11663_ _04011_ _04421_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__nor2_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _06121_ _06125_ _06124_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__a21bo_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10614_ _03645_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17170_ rbzero.traced_texa\[-1\] _09768_ _09769_ rbzero.wall_tracer.visualWallDist\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__a22o_1
X_14382_ _07117_ _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__or2_1
XFILLER_70_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11594_ _04242_ _04363_ _04372_ _04207_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__o211a_1
XFILLER_168_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16121_ _08765_ _08758_ vssd1 vssd1 vccd1 vccd1 _08766_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13333_ _06057_ _06067_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__nor2_1
X_10545_ _03609_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16052_ _08688_ _08683_ vssd1 vssd1 vccd1 vccd1 _08697_ sky130_fd_sc_hd__xnor2_1
XFILLER_115_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13264_ _05943_ _06000_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__xnor2_1
X_10476_ _03573_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15003_ rbzero.wall_tracer.stepDistX\[8\] _07579_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07672_ sky130_fd_sc_hd__mux2_1
X_12215_ _04960_ net16 net17 vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__a21o_1
XFILLER_123_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13195_ _05928_ _05901_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__or2_1
XFILLER_151_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19811_ _03134_ vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__clkbuf_1
X_12146_ net11 _04912_ _04914_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__o211ai_2
XFILLER_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03311_ clknet_0__03311_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03311_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_150_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19742_ rbzero.pov.spi_buffer\[45\] rbzero.pov.spi_buffer\[46\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03099_ sky130_fd_sc_hd__mux2_1
X_12077_ net7 _04848_ net3 net4 vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__and4b_1
X_16954_ _09342_ _09328_ _09456_ vssd1 vssd1 vccd1 vccd1 _09595_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15905_ _08509_ _08544_ vssd1 vssd1 vccd1 vccd1 _08550_ sky130_fd_sc_hd__xnor2_4
X_11028_ rbzero.tex_b0\[44\] rbzero.tex_b0\[43\] _03854_ vssd1 vssd1 vccd1 vccd1 _03863_
+ sky130_fd_sc_hd__mux2_1
X_19673_ rbzero.pov.spi_buffer\[12\] rbzero.pov.spi_buffer\[13\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03063_ sky130_fd_sc_hd__mux2_1
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16885_ _08705_ vssd1 vssd1 vccd1 vccd1 _09526_ sky130_fd_sc_hd__clkbuf_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18624_ _02319_ _02320_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__xor2_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _07958_ _08104_ vssd1 vssd1 vccd1 vccd1 _08481_ sky130_fd_sc_hd__nor2_1
XFILLER_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18555_ _02184_ _02196_ _02251_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a21o_1
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _08371_ _08411_ vssd1 vssd1 vccd1 vccd1 _08412_ sky130_fd_sc_hd__xor2_2
XFILLER_33_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12979_ _05710_ _05713_ _05715_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__or3_1
XFILLER_80_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17506_ _10071_ _09961_ vssd1 vssd1 vccd1 vccd1 _10072_ sky130_fd_sc_hd__nand2_1
XFILLER_61_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14718_ _07406_ _07432_ _07434_ _07454_ _05929_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__a32o_4
X_18486_ _02182_ _02183_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__and2_1
X_15698_ _08340_ _08341_ _08342_ vssd1 vssd1 vccd1 vccd1 _08343_ sky130_fd_sc_hd__and3_1
XFILLER_21_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17437_ _09709_ _09712_ vssd1 vssd1 vccd1 vccd1 _10004_ sky130_fd_sc_hd__nor2_1
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14649_ _07384_ _07385_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__or2_1
XANTENNA_16 _08094_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_38 net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ _09933_ _09934_ vssd1 vssd1 vccd1 vccd1 _09935_ sky130_fd_sc_hd__and2_1
XANTENNA_49 _08159_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19107_ rbzero.spi_registers.spi_buffer\[9\] rbzero.spi_registers.spi_buffer\[8\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__mux2_1
X_16319_ _08962_ _08963_ vssd1 vssd1 vccd1 vccd1 _08964_ sky130_fd_sc_hd__xnor2_1
XFILLER_203_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17299_ rbzero.wall_tracer.trackDistX\[-5\] _09870_ _05413_ vssd1 vssd1 vccd1 vccd1
+ _09871_ sky130_fd_sc_hd__mux2_1
XFILLER_174_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19038_ rbzero.pov.spi_buffer\[50\] rbzero.pov.ready_buffer\[50\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02651_ sky130_fd_sc_hd__mux2_1
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21000_ clknet_leaf_10_i_clk _00769_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20715_ clknet_leaf_47_i_clk _00016_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_178_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20646_ clknet_leaf_62_i_clk _00430_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_177_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20577_ _02721_ _03448_ _03449_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__and3_1
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10330_ rbzero.tex_r1\[53\] rbzero.tex_r1\[54\] _03494_ vssd1 vssd1 vccd1 vccd1 _03495_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12000_ rbzero.tex_b1\[55\] rbzero.tex_b1\[54\] _04250_ vssd1 vssd1 vccd1 vccd1 _04775_
+ sky130_fd_sc_hd__mux2_1
XFILLER_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21129_ clknet_leaf_4_i_clk _00898_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13951_ _06675_ _06672_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__nor2_1
XFILLER_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12902_ _05562_ _05566_ _05601_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__and3_1
X_16670_ _09149_ _09151_ vssd1 vssd1 vccd1 vccd1 _09313_ sky130_fd_sc_hd__and2b_1
X_13882_ _06568_ _06586_ _06587_ _06618_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__a31o_1
XFILLER_189_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15621_ _07988_ vssd1 vssd1 vccd1 vccd1 _08266_ sky130_fd_sc_hd__clkinv_2
XFILLER_62_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12833_ rbzero.wall_tracer.rcp_sel\[2\] vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__inv_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _01737_ _10238_ _09294_ _09977_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__or4_1
XFILLER_61_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _05510_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__clkbuf_1
X_15552_ _07549_ _07552_ _07555_ vssd1 vssd1 vccd1 vccd1 _08197_ sky130_fd_sc_hd__and3_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11715_ rbzero.debug_overlay.facingX\[-6\] _04475_ _04458_ rbzero.debug_overlay.facingX\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__a22o_1
X_14503_ _06239_ _07071_ _07238_ _07239_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__or4bb_1
X_18271_ _01756_ _01970_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__xnor2_4
XFILLER_188_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15483_ _08125_ vssd1 vssd1 vccd1 vccd1 _08128_ sky130_fd_sc_hd__clkbuf_4
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ rbzero.debug_overlay.facingX\[0\] rbzero.wall_tracer.rayAddendX\[8\] vssd1
+ vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__nand2_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17222_ _09800_ _09801_ vssd1 vssd1 vccd1 vccd1 _09802_ sky130_fd_sc_hd__xnor2_1
X_11646_ gpout0.hpos\[4\] _04024_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__nor2_1
X_14434_ _06153_ _06705_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__and2_1
XFILLER_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput14 i_gpout2_sel[0] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_6
XFILLER_168_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17153_ rbzero.row_render.texu\[3\] _09766_ _07728_ net511 vssd1 vssd1 vccd1 vccd1
+ _00542_ sky130_fd_sc_hd__a22o_1
Xinput25 i_gpout3_sel[5] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__buf_6
X_14365_ _05793_ _07101_ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__nor2_1
Xinput36 i_gpout5_sel[4] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_4
X_11577_ _04341_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__buf_6
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput47 i_tex_in[1] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_4
X_16104_ _08745_ _08746_ _08748_ vssd1 vssd1 vccd1 vccd1 _08749_ sky130_fd_sc_hd__a21boi_2
X_13316_ _05939_ _06052_ _05922_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__or3b_4
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10528_ _03600_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__clkbuf_1
X_17084_ _09538_ _09578_ _09723_ vssd1 vssd1 vccd1 vccd1 _09724_ sky130_fd_sc_hd__a21boi_2
XFILLER_122_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14296_ _06703_ _06841_ _07032_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__a21oi_2
XFILLER_109_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13247_ _05945_ _05949_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__and2_2
X_16035_ _08631_ _08675_ _08678_ _08679_ vssd1 vssd1 vccd1 vccd1 _08680_ sky130_fd_sc_hd__o22a_1
X_10459_ _03564_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13178_ _05880_ _05882_ _05811_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__mux2_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12129_ _04871_ _04881_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__or3_2
X_17986_ _01580_ _01590_ _01588_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__a21o_1
XFILLER_69_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19725_ rbzero.pov.spi_buffer\[37\] rbzero.pov.spi_buffer\[38\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03090_ sky130_fd_sc_hd__mux2_1
XFILLER_81_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16937_ _09575_ _09577_ vssd1 vssd1 vccd1 vccd1 _09578_ sky130_fd_sc_hd__xnor2_1
XFILLER_78_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19656_ rbzero.pov.spi_buffer\[4\] rbzero.pov.spi_buffer\[5\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03054_ sky130_fd_sc_hd__mux2_1
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16868_ _09363_ _09371_ _09508_ vssd1 vssd1 vccd1 vccd1 _09509_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18607_ _02301_ _02302_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__and2_1
XFILLER_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15819_ _08440_ _08463_ vssd1 vssd1 vccd1 vccd1 _08464_ sky130_fd_sc_hd__nand2_1
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20263__281 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__inv_2
X_16799_ _09439_ _09440_ vssd1 vssd1 vccd1 vccd1 _09441_ sky130_fd_sc_hd__xor2_2
XFILLER_92_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18538_ _02141_ _02160_ _02140_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__a21bo_1
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18469_ _10094_ _09350_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__nor2_1
XFILLER_21_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20500_ _03395_ _03396_ _03397_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__and3_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21480_ net401 _01249_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_53_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20431_ _03338_ _03339_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__nand2_1
XFILLER_53_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20346__356 clknet_1_0__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__inv_2
XFILLER_21_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11500_ _04277_ _04278_ _04279_ _04226_ _04210_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__o221a_1
XFILLER_196_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12480_ _05214_ rbzero.wall_tracer.trackDistX\[10\] _05224_ rbzero.wall_tracer.trackDistY\[4\]
+ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__a221o_1
Xclkbuf_1_0__f__03314_ clknet_0__03314_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03314_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _04128_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__buf_4
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20629_ clknet_leaf_14_i_clk _00413_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14150_ _06862_ _06869_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__xnor2_2
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11362_ _04097_ _04114_ _04117_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__nor3_4
X_20091__126 clknet_1_0__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__inv_2
X_13101_ _05836_ _05837_ _05807_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__mux2_1
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10313_ rbzero.tex_r1\[61\] rbzero.tex_r1\[62\] _03483_ vssd1 vssd1 vccd1 vccd1 _03486_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_1_0_i_clk clknet_1_0_1_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_164_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14081_ _06737_ _06817_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__xnor2_2
X_11293_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] vssd1 vssd1
+ vccd1 vccd1 _04073_ sky130_fd_sc_hd__nand2_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _05691_ _05673_ _05683_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__or4_1
XFILLER_106_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17840_ _10281_ _10283_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__nor2_1
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17771_ _08157_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__clkbuf_4
X_14983_ rbzero.wall_tracer.stepDistX\[-2\] _07650_ vssd1 vssd1 vccd1 vccd1 _07662_
+ sky130_fd_sc_hd__nor2_1
XFILLER_75_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19510_ _07679_ _02978_ _02979_ _02988_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__a31o_1
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16722_ _09244_ _09248_ vssd1 vssd1 vccd1 vccd1 _09364_ sky130_fd_sc_hd__nand2_1
X_13934_ _06607_ _06610_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__xor2_4
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19441_ _02904_ rbzero.wall_tracer.rayAddendY\[3\] vssd1 vssd1 vccd1 vccd1 _02924_
+ sky130_fd_sc_hd__nor2_1
X_16653_ _08239_ _09135_ _09294_ _09295_ vssd1 vssd1 vccd1 vccd1 _09296_ sky130_fd_sc_hd__o31ai_1
X_13865_ _06425_ _06555_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__nand2_2
XFILLER_62_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__03041_ _03041_ vssd1 vssd1 vccd1 vccd1 clknet_0__03041_ sky130_fd_sc_hd__clkbuf_16
X_15604_ _08206_ _08248_ vssd1 vssd1 vccd1 vccd1 _08249_ sky130_fd_sc_hd__xnor2_4
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19372_ rbzero.debug_overlay.vplaneY\[-2\] rbzero.wall_tracer.rayAddendY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__or2_1
X_12816_ _05548_ _05552_ _05554_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__o21ai_1
XFILLER_188_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16584_ _09225_ _09226_ vssd1 vssd1 vccd1 vccd1 _09227_ sky130_fd_sc_hd__nand2_1
X_13796_ _05855_ _05877_ _06061_ _06078_ _06532_ vssd1 vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__a41o_1
XFILLER_62_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18323_ _02016_ _02022_ rbzero.wall_tracer.trackDistX\[7\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00596_ sky130_fd_sc_hd__o2bb2a_1
X_15535_ _07989_ vssd1 vssd1 vccd1 vccd1 _08180_ sky130_fd_sc_hd__buf_4
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _05454_ _05456_ _05491_ _05494_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a31o_4
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _08257_ _08242_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__or4_1
X_15466_ _08109_ vssd1 vssd1 vccd1 vccd1 _08111_ sky130_fd_sc_hd__buf_4
X_12678_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__nand2_1
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17205_ rbzero.wall_tracer.mapX\[8\] _05525_ vssd1 vssd1 vccd1 vccd1 _09788_ sky130_fd_sc_hd__xor2_1
X_11629_ _04402_ _04404_ _04407_ _04306_ _04241_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a221o_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14417_ _07146_ _07153_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__and2_1
XFILLER_204_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18185_ _10271_ _01766_ _01884_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__or3b_1
XFILLER_200_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15397_ _08041_ vssd1 vssd1 vccd1 vccd1 _08042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_11_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17136_ _07855_ vssd1 vssd1 vccd1 vccd1 _09764_ sky130_fd_sc_hd__buf_2
XFILLER_190_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14348_ _07059_ _07083_ vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__or2_1
XFILLER_116_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17067_ _09704_ _09705_ _09706_ vssd1 vssd1 vccd1 vccd1 _09707_ sky130_fd_sc_hd__a21bo_2
X_14279_ _06666_ _06760_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__nor2_1
XFILLER_98_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16018_ _08658_ _08662_ vssd1 vssd1 vccd1 vccd1 _08663_ sky130_fd_sc_hd__xor2_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _10292_ _01671_ _01549_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__a21o_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19708_ _03047_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__buf_4
X_20980_ clknet_leaf_13_i_clk _00749_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03308_ _03308_ vssd1 vssd1 vccd1 vccd1 clknet_0__03308_ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21601_ net142 _01370_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21532_ net453 _01301_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21463_ net384 _01232_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20414_ rbzero.traced_texa\[-12\] rbzero.texV\[-12\] vssd1 vssd1 vccd1 vccd1 _03326_
+ sky130_fd_sc_hd__or2_1
XFILLER_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21394_ net315 _01163_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19639__89 clknet_1_0__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__inv_2
XFILLER_108_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ rbzero.tex_b1\[14\] _04338_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__and2_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10931_ _03812_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10862_ _03776_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__clkbuf_1
X_13650_ _06381_ _06386_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__and2b_1
XFILLER_72_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12601_ _05352_ _05354_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__and2_1
X_13581_ _06288_ _06317_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__nor2_1
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _03717_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__clkbuf_4
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12532_ rbzero.debug_overlay.facingY\[0\] rbzero.wall_tracer.rayAddendY\[8\] vssd1
+ vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__or2_1
X_15320_ _05196_ rbzero.wall_tracer.stepDistX\[-6\] vssd1 vssd1 vccd1 vccd1 _07965_
+ sky130_fd_sc_hd__nor2_2
XFILLER_157_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12463_ rbzero.wall_tracer.trackDistX\[7\] vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__inv_2
X_15251_ _07895_ _07595_ _07896_ _07642_ vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__o211a_1
XFILLER_138_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_81 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_81/HI o_rgb[11] sky130_fd_sc_hd__conb_1
X_11414_ rbzero.row_render.size\[1\] _04192_ _04193_ _04148_ vssd1 vssd1 vccd1 vccd1
+ _04194_ sky130_fd_sc_hd__a211o_1
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14202_ _06926_ _06935_ _06938_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__a21boi_1
Xtop_ew_algofoogle_92 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_92/HI zeros[2] sky130_fd_sc_hd__conb_1
XFILLER_138_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15182_ _07820_ _04462_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1
+ _07836_ sky130_fd_sc_hd__or3b_1
X_12394_ net46 _05144_ _05139_ _04323_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a22o_1
XFILLER_184_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14133_ _06863_ _06868_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__or2b_1
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ _04089_ _04114_ _04124_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__or3b_4
XFILLER_193_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19990_ rbzero.pov.ready_buffer\[16\] _03246_ _03248_ rbzero.debug_overlay.vplaneX\[-4\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_94_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_141_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14064_ _06666_ _06663_ _06712_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__o21ai_1
X_18941_ rbzero.pov.spi_buffer\[4\] rbzero.pov.ready_buffer\[4\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02600_ sky130_fd_sc_hd__mux2_1
X_11276_ rbzero.texV\[8\] _04054_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__a21boi_1
XFILLER_165_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13015_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__buf_4
XFILLER_121_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18872_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.stepDistY\[10\] vssd1
+ vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__nand2_1
X_17823_ _09117_ _10266_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__nor2_1
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20329__340 clknet_1_0__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__inv_2
Xhold3 rbzero.wall_tracer.texu\[3\] vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17754_ _09249_ _09480_ _09484_ _09096_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__o22a_1
XFILLER_82_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14966_ rbzero.wall_tracer.stepDistX\[-10\] _07484_ _07650_ vssd1 vssd1 vccd1 vccd1
+ _07653_ sky130_fd_sc_hd__mux2_1
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16705_ _09345_ _09346_ vssd1 vssd1 vccd1 vccd1 _09347_ sky130_fd_sc_hd__nor2_1
X_13917_ _06616_ _06595_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__nand2_1
X_17685_ _09126_ _10248_ _10100_ _10249_ vssd1 vssd1 vccd1 vccd1 _10250_ sky130_fd_sc_hd__o31a_1
XFILLER_75_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14897_ rbzero.wall_tracer.trackDistY\[-8\] rbzero.wall_tracer.trackDistX\[-8\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__mux2_1
XFILLER_207_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_19424_ _02893_ _02896_ _02907_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a21oi_1
XFILLER_207_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16636_ _05209_ rbzero.wall_tracer.stepDistX\[5\] vssd1 vssd1 vccd1 vccd1 _09279_
+ sky130_fd_sc_hd__nand2_2
X_13848_ _06583_ _06584_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__nor2_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19355_ _02843_ _02844_ _07703_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__a21oi_1
XFILLER_62_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16567_ _09090_ _09112_ _09110_ vssd1 vssd1 vccd1 vccd1 _09210_ sky130_fd_sc_hd__a21o_1
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13779_ _05855_ _06153_ _06501_ _06502_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__a22o_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18306_ _01928_ _02005_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15518_ _08162_ _08159_ _08160_ _08151_ vssd1 vssd1 vccd1 vccd1 _08163_ sky130_fd_sc_hd__o22a_1
XFILLER_148_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19286_ rbzero.spi_registers.spi_buffer\[5\] rbzero.spi_registers.new_leak\[5\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__mux2_1
XFILLER_203_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16498_ _08977_ _08978_ vssd1 vssd1 vccd1 vccd1 _09142_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_47_i_clk clknet_3_4_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18237_ _09526_ _09703_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__nand2_1
X_20375__382 clknet_1_0__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__inv_2
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15449_ _08093_ rbzero.debug_overlay.playerX\[-1\] _05496_ vssd1 vssd1 vccd1 vccd1
+ _08094_ sky130_fd_sc_hd__mux2_1
XFILLER_50_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18168_ _09674_ _09693_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__nor2_1
X_20074__110 clknet_1_0__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__inv_2
XFILLER_11_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17119_ _09755_ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18099_ _01684_ _01685_ _01785_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__a21o_1
XFILLER_143_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20061_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__buf_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20963_ clknet_leaf_5_i_clk _00732_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20894_ clknet_leaf_86_i_clk _00663_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21515_ net436 _01284_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21446_ net367 _01215_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21377_ net298 _01146_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11130_ rbzero.map_rom.f4 vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__clkinv_2
XFILLER_107_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11061_ _03880_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_131_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ _07547_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__clkbuf_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _07485_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__clkbuf_1
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11963_ _04738_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__inv_2
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _06396_ _06413_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__xor2_1
X_10914_ _03803_ vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__clkbuf_1
X_17470_ _10028_ _10035_ rbzero.wall_tracer.trackDistX\[0\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00589_ sky130_fd_sc_hd__o2bb2a_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14682_ _07107_ _07413_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__nand2_2
X_11894_ _04667_ _04668_ _04669_ _04379_ _04332_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__o221a_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16421_ _09064_ _09065_ vssd1 vssd1 vccd1 vccd1 _09066_ sky130_fd_sc_hd__or2b_1
X_13633_ _06351_ _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__nor2_1
X_10845_ _03767_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19140_ _04890_ _04315_ _02703_ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__nor4_4
X_16352_ _08281_ _08296_ _08996_ vssd1 vssd1 vccd1 vccd1 _08997_ sky130_fd_sc_hd__a21oi_4
X_10776_ _03731_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13564_ _06284_ _06300_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15303_ _07946_ _07947_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__nand2_1
X_19071_ rbzero.pov.spi_buffer\[66\] rbzero.pov.ready_buffer\[66\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02668_ sky130_fd_sc_hd__mux2_1
X_12515_ rbzero.wall_tracer.trackDistY\[-3\] _05267_ _05263_ rbzero.wall_tracer.trackDistY\[-4\]
+ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__o221a_1
X_16283_ _08924_ _08926_ vssd1 vssd1 vccd1 vccd1 _08928_ sky130_fd_sc_hd__nand2_1
XFILLER_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13495_ _06230_ _06196_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__and2b_1
XFILLER_201_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18022_ _01717_ _01619_ _01723_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a21oi_1
XFILLER_173_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15234_ _07882_ _07883_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__nor2_1
X_12446_ net71 rbzero.wall_tracer.state\[2\] _05190_ vssd1 vssd1 vccd1 vccd1 _05202_
+ sky130_fd_sc_hd__and3_1
XFILLER_139_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12377_ _05141_ _05143_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__nor2_1
XFILLER_125_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15165_ _07785_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__buf_2
XFILLER_5_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11328_ _04053_ _04056_ _04107_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__o21a_1
X_14116_ _06692_ _06852_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__and2_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15096_ rbzero.wall_tracer.rayAddendX\[0\] _00013_ _07747_ _07755_ vssd1 vssd1 vccd1
+ vccd1 _00496_ sky130_fd_sc_hd__o22a_1
XFILLER_10_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19973_ rbzero.pov.ready_buffer\[24\] _03247_ _03249_ rbzero.debug_overlay.facingY\[-7\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__a221o_1
XFILLER_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18924_ rbzero.spi_registers.spi_counter\[5\] rbzero.spi_registers.spi_counter\[4\]
+ _02583_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__and3_1
X_14047_ _06768_ _06783_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__xnor2_1
X_11259_ rbzero.wall_tracer.state\[10\] _04038_ _04039_ vssd1 vssd1 vccd1 vccd1 _00014_
+ sky130_fd_sc_hd__o21a_1
XFILLER_141_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18855_ rbzero.wall_tracer.trackDistY\[8\] rbzero.wall_tracer.stepDistY\[8\] vssd1
+ vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__nor2_1
XFILLER_94_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17806_ _01507_ _01509_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__xor2_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18786_ _02464_ _02398_ _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__and3_1
XFILLER_36_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15998_ _07601_ _04014_ _07990_ _07936_ vssd1 vssd1 vccd1 vccd1 _08643_ sky130_fd_sc_hd__and4_1
XFILLER_95_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17737_ _10186_ _10288_ _01440_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__a21o_1
X_14949_ _07621_ _07640_ _07641_ _07642_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__o211a_1
XFILLER_78_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17668_ _10197_ _10232_ vssd1 vssd1 vccd1 vccd1 _10233_ sky130_fd_sc_hd__xnor2_1
XFILLER_39_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20106__139 clknet_1_1__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__inv_2
X_19407_ rbzero.wall_tracer.rayAddendY\[0\] _00013_ _02892_ vssd1 vssd1 vccd1 vccd1
+ _00810_ sky130_fd_sc_hd__o21a_1
X_16619_ _09251_ _09261_ vssd1 vssd1 vccd1 vccd1 _09262_ sky130_fd_sc_hd__xnor2_1
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17599_ _10037_ _10038_ _10164_ vssd1 vssd1 vccd1 vccd1 _10165_ sky130_fd_sc_hd__and3_1
XFILLER_204_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19338_ rbzero.debug_overlay.vplaneY\[-8\] rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__nand2_1
XFILLER_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19269_ _02788_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21300_ net221 _01069_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21231_ clknet_leaf_17_i_clk _01000_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_117_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21162_ clknet_leaf_86_i_clk _00931_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21093_ net183 _00862_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19617__70 clknet_1_0__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__inv_2
X_20044_ _04886_ _03278_ _04887_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__a21o_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19632__84 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__inv_2
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_0_0_i_clk clknet_2_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_113_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20946_ clknet_leaf_4_i_clk _00715_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ clknet_leaf_96_i_clk _00646_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10630_ _03654_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10561_ rbzero.tex_r0\[10\] rbzero.tex_r0\[9\] _03613_ vssd1 vssd1 vccd1 vccd1 _03618_
+ sky130_fd_sc_hd__mux2_1
X_12300_ _05066_ _05067_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__or3b_2
XFILLER_194_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13280_ _06015_ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__or2_1
X_10492_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _03580_ vssd1 vssd1 vccd1 vccd1 _03582_
+ sky130_fd_sc_hd__mux2_1
XFILLER_154_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ net125 _04960_ _04966_ net17 net16 vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a2111o_2
X_21429_ net350 _01198_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12162_ _04317_ _04931_ _04932_ net9 net11 vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__o221a_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11113_ _03907_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_111_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12093_ net5 net4 vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__nor2_1
X_20211__234 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__inv_2
X_16970_ rbzero.wall_tracer.visualWallDist\[11\] _04015_ vssd1 vssd1 vccd1 vccd1 _09610_
+ sky130_fd_sc_hd__nand2_1
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15921_ _08557_ _08563_ _08565_ vssd1 vssd1 vccd1 vccd1 _08566_ sky130_fd_sc_hd__a21o_1
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11044_ _03871_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_103_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18640_ _09284_ _09287_ _08151_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__a21o_1
XFILLER_76_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _08097_ _08491_ vssd1 vssd1 vccd1 vccd1 _08497_ sky130_fd_sc_hd__nor2_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14803_ _07473_ _07499_ _07532_ _07527_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__o211a_1
XFILLER_188_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ _02259_ _02267_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__xor2_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _08135_ _08427_ _08422_ vssd1 vssd1 vccd1 vccd1 _08428_ sky130_fd_sc_hd__o21ai_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ _05703_ _05722_ _05727_ _05731_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a211o_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ _10050_ _10087_ vssd1 vssd1 vccd1 vccd1 _10088_ sky130_fd_sc_hd__xnor2_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14734_ _07378_ _07413_ _07415_ vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__a21o_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ rbzero.tex_b0\[47\] _04347_ _04348_ _04217_ vssd1 vssd1 vccd1 vccd1 _04722_
+ sky130_fd_sc_hd__a31o_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ _09726_ _09728_ vssd1 vssd1 vccd1 vccd1 _10020_ sky130_fd_sc_hd__nor2_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _07386_ _07401_ _05779_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__mux2_1
X_11877_ rbzero.tex_g1\[25\] rbzero.tex_g1\[24\] _04336_ vssd1 vssd1 vccd1 vccd1 _04654_
+ sky130_fd_sc_hd__mux2_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16404_ _09047_ _09048_ vssd1 vssd1 vccd1 vccd1 _09049_ sky130_fd_sc_hd__xnor2_4
X_13616_ _06319_ _06316_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__or2b_1
X_17384_ _09938_ _09950_ vssd1 vssd1 vccd1 vccd1 _09951_ sky130_fd_sc_hd__xnor2_1
X_10828_ _03758_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__clkbuf_1
X_14596_ _07216_ _07331_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__nor2_1
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19123_ _02696_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__clkbuf_1
X_16335_ _08230_ rbzero.wall_tracer.stepDistY\[6\] vssd1 vssd1 vccd1 vccd1 _08980_
+ sky130_fd_sc_hd__nand2_1
XFILLER_119_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13547_ _06136_ _06137_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__xor2_1
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10759_ _03722_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19054_ rbzero.pov.spi_buffer\[58\] rbzero.pov.ready_buffer\[58\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02659_ sky130_fd_sc_hd__mux2_1
X_16266_ _08853_ _08910_ vssd1 vssd1 vccd1 vccd1 _08911_ sky130_fd_sc_hd__nor2_1
XFILLER_195_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13478_ _05990_ _06134_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__nor2_1
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18005_ _01582_ _01706_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__xnor2_1
X_15217_ _07845_ _07864_ vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__nor2_1
X_12429_ _05191_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__clkbuf_1
X_16197_ _08840_ _08841_ vssd1 vssd1 vccd1 vccd1 _08842_ sky130_fd_sc_hd__nor2_1
XFILLER_127_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15148_ _07802_ _07803_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__nor2_1
XFILLER_141_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15079_ rbzero.wall_tracer.rayAddendX\[-1\] _07706_ _07739_ _07703_ vssd1 vssd1 vccd1
+ vccd1 _07740_ sky130_fd_sc_hd__a22o_1
X_19956_ rbzero.pov.ready_buffer\[36\] _03240_ _03243_ rbzero.debug_overlay.facingX\[-6\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__o221a_1
XFILLER_113_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20186__211 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__inv_2
X_18907_ _02574_ _02575_ _02576_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__and3_1
XFILLER_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19887_ rbzero.debug_overlay.playerY\[-9\] vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__inv_2
XFILLER_56_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18838_ rbzero.wall_tracer.trackDistY\[5\] _02515_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02516_ sky130_fd_sc_hd__mux2_1
XFILLER_67_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18769_ rbzero.wall_tracer.trackDistY\[-4\] _02455_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02456_ sky130_fd_sc_hd__mux2_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20800_ clknet_leaf_44_i_clk _00569_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.wall\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20731_ clknet_leaf_68_i_clk _00500_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20662_ clknet_leaf_63_i_clk _00446_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20593_ _07679_ _02832_ _03459_ _07855_ rbzero.wall_tracer.rayAddendY\[-8\] vssd1
+ vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__a32o_1
XFILLER_192_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21214_ clknet_leaf_22_i_clk _00983_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21145_ clknet_leaf_97_i_clk _00914_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21076_ net166 _00845_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20027_ _04892_ _04992_ _04883_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ rbzero.tex_g0\[47\] _04135_ _04136_ _04126_ vssd1 vssd1 vccd1 vccd1 _04578_
+ sky130_fd_sc_hd__a31o_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12780_ _05524_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__clkbuf_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ rbzero.debug_overlay.playerX\[-7\] _04455_ _04458_ rbzero.debug_overlay.playerX\[-9\]
+ _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__a221o_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20929_ clknet_leaf_26_i_clk _00698_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _06153_ _07072_ _07186_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a21o_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ gpout0.hpos\[7\] _04414_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__nor2_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13401_ _06136_ _06137_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__or2b_1
X_10613_ rbzero.tex_g1\[48\] rbzero.tex_g1\[49\] _03635_ vssd1 vssd1 vccd1 vccd1 _03645_
+ sky130_fd_sc_hd__mux2_1
X_11593_ _04254_ _04366_ _04370_ _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__a211o_1
X_14381_ _06696_ _06760_ _07116_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__o21ba_1
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16120_ _08759_ _08756_ vssd1 vssd1 vccd1 vccd1 _08765_ sky130_fd_sc_hd__and2b_1
XFILLER_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10544_ rbzero.tex_r0\[18\] rbzero.tex_r0\[17\] _03602_ vssd1 vssd1 vccd1 vccd1 _03609_
+ sky130_fd_sc_hd__mux2_1
X_13332_ _06058_ _06063_ _06064_ _06068_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16051_ _08638_ _08651_ vssd1 vssd1 vccd1 vccd1 _08696_ sky130_fd_sc_hd__xnor2_1
X_10475_ rbzero.tex_r0\[51\] rbzero.tex_r0\[50\] _03569_ vssd1 vssd1 vccd1 vccd1 _03573_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13263_ _05998_ _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__nor2_1
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15002_ _07671_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12214_ net18 net19 _04983_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__and3b_1
XFILLER_124_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13194_ _05826_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__buf_2
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ _04910_ net66 _04915_ net12 vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__a211o_1
X_19810_ rbzero.pov.sclk_buffer\[1\] rbzero.pov.sclk_buffer\[0\] _05189_ vssd1 vssd1
+ vccd1 vccd1 _03134_ sky130_fd_sc_hd__mux2_1
XFILLER_151_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03310_ clknet_0__03310_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03310_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12076_ _04840_ net64 _04846_ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__a211o_1
XFILLER_173_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16953_ _09592_ _09593_ vssd1 vssd1 vccd1 vccd1 _09594_ sky130_fd_sc_hd__nor2_4
X_19741_ _03098_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__clkbuf_1
X_15904_ _08547_ _08548_ vssd1 vssd1 vccd1 vccd1 _08549_ sky130_fd_sc_hd__nor2_4
X_11027_ _03862_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__clkbuf_1
X_19672_ _03062_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__clkbuf_1
X_16884_ _08705_ _08059_ _09524_ vssd1 vssd1 vccd1 vccd1 _09525_ sky130_fd_sc_hd__or3_1
XFILLER_37_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18623_ _02229_ _02231_ _02230_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__a21boi_1
X_20406__7 clknet_1_1__leaf__03037_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__inv_2
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _07913_ _07967_ _08022_ _07923_ vssd1 vssd1 vccd1 vccd1 _08480_ sky130_fd_sc_hd__o22ai_1
XFILLER_65_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19611__65 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__inv_2
X_18554_ _02193_ _02195_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__nor2_1
X_15766_ _08400_ _08409_ _08410_ vssd1 vssd1 vccd1 vccd1 _08411_ sky130_fd_sc_hd__a21oi_2
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12978_ _05584_ _05714_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__xor2_2
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17505_ _09663_ _09959_ vssd1 vssd1 vccd1 vccd1 _10071_ sky130_fd_sc_hd__or2_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14717_ _07439_ _07444_ _07449_ _07453_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__nand4_1
X_18485_ _02171_ _02181_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__or2_1
X_11929_ rbzero.tex_b0\[56\] _04338_ _04225_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__a21o_1
X_15697_ _08097_ _08022_ vssd1 vssd1 vccd1 vccd1 _08342_ sky130_fd_sc_hd__nor2_1
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17436_ _09994_ _10002_ vssd1 vssd1 vccd1 vccd1 _10003_ sky130_fd_sc_hd__xnor2_1
X_14648_ _05893_ _07365_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__and2_1
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _08283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17367_ _09931_ _09932_ vssd1 vssd1 vccd1 vccd1 _09934_ sky130_fd_sc_hd__nand2_1
XANTENNA_39 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ _07285_ _07293_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__nand2_1
XFILLER_158_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19106_ _02686_ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__clkbuf_1
X_16318_ _07913_ _08264_ vssd1 vssd1 vccd1 vccd1 _08963_ sky130_fd_sc_hd__and2b_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17298_ _09863_ _09867_ _09868_ _09869_ vssd1 vssd1 vccd1 vccd1 _09870_ sky130_fd_sc_hd__o31ai_1
X_19037_ _02650_ vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__clkbuf_1
X_16249_ _08877_ _08878_ vssd1 vssd1 vccd1 vccd1 _08894_ sky130_fd_sc_hd__or2b_1
XFILLER_134_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19939_ _02820_ _03232_ _03197_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__o21a_1
XFILLER_102_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20240__260 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__inv_2
XFILLER_54_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20714_ clknet_leaf_71_i_clk _00005_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20645_ clknet_leaf_62_i_clk _00429_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20576_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__or2_1
XFILLER_178_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20158__187 clknet_1_1__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__inv_2
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21128_ clknet_leaf_94_i_clk _00897_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13950_ _06685_ _06686_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__nand2_1
X_21059_ clknet_leaf_0_i_clk _00828_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12901_ _05632_ _05634_ _05636_ _05637_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__or4b_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13881_ _06591_ _06589_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__and2b_1
XFILLER_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15620_ _08263_ _08264_ vssd1 vssd1 vccd1 vccd1 _08265_ sky130_fd_sc_hd__and2_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20323__335 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__inv_2
XFILLER_185_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12832_ _04031_ _05372_ _05568_ _04001_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__a211o_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _07894_ _05459_ _08195_ _05193_ vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__a211o_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12763_ rbzero.map_rom.f2 _05509_ _05414_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__mux2_1
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _06002_ _06770_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__nand2_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _01969_ _10110_ _01879_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__mux2_2
XFILLER_187_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11714_ rbzero.debug_overlay.facingX\[-3\] _04463_ _04466_ rbzero.debug_overlay.facingX\[-8\]
+ _04481_ vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__a221o_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15482_ _08126_ vssd1 vssd1 vccd1 vccd1 _08127_ sky130_fd_sc_hd__inv_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12694_ _05418_ _05439_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__nand3b_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ rbzero.wall_tracer.mapX\[11\] _05525_ vssd1 vssd1 vccd1 vccd1 _09801_ sky130_fd_sc_hd__xnor2_1
X_14433_ _07142_ _07169_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__or2_1
X_11645_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__inv_2
XFILLER_168_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17152_ rbzero.row_render.texu\[2\] _09766_ _07728_ rbzero.wall_tracer.texu\[2\]
+ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__a22o_1
Xinput15 i_gpout2_sel[1] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_6
X_14364_ _07099_ _07100_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__or2_1
XFILLER_161_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11576_ _04232_ _04333_ _04340_ _04354_ _04244_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__o311a_1
Xinput26 i_gpout4_sel[0] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_4
XFILLER_11_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 i_gpout5_sel[5] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_4
Xinput48 i_tex_in[2] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_4
XFILLER_156_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16103_ _07964_ _08674_ _08747_ vssd1 vssd1 vccd1 vccd1 _08748_ sky130_fd_sc_hd__or3_1
X_13315_ _05973_ _05961_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__or2_1
X_10527_ rbzero.tex_r0\[26\] rbzero.tex_r0\[25\] _03591_ vssd1 vssd1 vccd1 vccd1 _03600_
+ sky130_fd_sc_hd__mux2_1
X_17083_ _09575_ _09577_ vssd1 vssd1 vccd1 vccd1 _09723_ sky130_fd_sc_hd__or2b_1
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14295_ _06818_ _06840_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__nor2_1
XFILLER_155_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16034_ _08008_ _08104_ vssd1 vssd1 vccd1 vccd1 _08679_ sky130_fd_sc_hd__or2_1
X_10458_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _03558_ vssd1 vssd1 vccd1 vccd1 _03564_
+ sky130_fd_sc_hd__mux2_1
X_13246_ _05961_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__buf_2
XFILLER_108_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10389_ _03525_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__clkbuf_1
X_13177_ _05902_ _05879_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__or2_1
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12128_ net7 _04882_ _04894_ _04899_ _04837_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__a32o_2
X_17985_ _01575_ _01607_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__or2_1
XFILLER_42_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12059_ _03474_ _04815_ _04005_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__o21ai_1
X_16936_ _09415_ _09441_ _09576_ vssd1 vssd1 vccd1 vccd1 _09577_ sky130_fd_sc_hd__a21o_1
X_19724_ _03089_ vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16867_ _09244_ _09248_ _09370_ vssd1 vssd1 vccd1 vccd1 _09508_ sky130_fd_sc_hd__a21oi_1
X_19655_ _03053_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18606_ _02301_ _02302_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__nor2_1
X_15818_ _08460_ _08461_ _08462_ vssd1 vssd1 vccd1 vccd1 _08463_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16798_ _09297_ _09299_ vssd1 vssd1 vccd1 vccd1 _09440_ sky130_fd_sc_hd__and2_1
XFILLER_129_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20298__312 clknet_1_1__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__inv_2
X_18537_ _02228_ _02234_ rbzero.wall_tracer.trackDistX\[9\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00598_ sky130_fd_sc_hd__o2bb2a_1
X_15749_ _08316_ _08314_ vssd1 vssd1 vccd1 vccd1 _08394_ sky130_fd_sc_hd__nand2_1
XFILLER_61_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18468_ _02038_ _02053_ _02165_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__a21bo_1
XFILLER_34_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17419_ _09975_ _09985_ vssd1 vssd1 vccd1 vccd1 _09986_ sky130_fd_sc_hd__xor2_2
XFILLER_166_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18399_ _02096_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__and2b_1
XFILLER_20_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20430_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 _03339_
+ sky130_fd_sc_hd__nand2_1
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20164__191 clknet_1_0__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__inv_2
XFILLER_58_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__03313_ clknet_0__03313_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03313_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ _04209_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__buf_4
X_20628_ clknet_leaf_24_i_clk _00412_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapX\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_193_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11361_ _04093_ _04114_ _04122_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__nor3_2
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20559_ _09763_ _09194_ rbzero.traced_texVinit\[3\] _09762_ vssd1 vssd1 vccd1 vccd1
+ _01411_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10312_ _03485_ vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__clkbuf_1
X_13100_ _05642_ _05645_ _05796_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__mux2_1
XFILLER_125_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14080_ _06798_ _06816_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__xnor2_2
X_11292_ rbzero.traced_texVinit\[4\] rbzero.spi_registers.vshift\[1\] vssd1 vssd1
+ vccd1 vccd1 _04072_ sky130_fd_sc_hd__or2_1
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13031_ _05642_ _05744_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__nand2_1
XFILLER_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17770_ _05198_ _08445_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__nand2_2
X_14982_ _07661_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__clkbuf_1
X_16721_ _09226_ _09228_ _09225_ vssd1 vssd1 vccd1 vccd1 _09363_ sky130_fd_sc_hd__a21bo_1
X_13933_ _06666_ _06668_ _06669_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__or3_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19440_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__and2_1
XFILLER_74_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16652_ _09133_ _09134_ vssd1 vssd1 vccd1 vccd1 _09295_ sky130_fd_sc_hd__or2_1
X_13864_ _06559_ _06378_ _06558_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__nand3_1
XFILLER_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__03040_ _03040_ vssd1 vssd1 vccd1 vccd1 clknet_0__03040_ sky130_fd_sc_hd__clkbuf_16
X_15603_ _08241_ _08247_ vssd1 vssd1 vccd1 vccd1 _08248_ sky130_fd_sc_hd__xor2_4
XFILLER_90_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19371_ _02859_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__clkbuf_1
X_12815_ rbzero.wall_tracer.mapY\[10\] _05404_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__xor2_1
X_16583_ _08823_ _08159_ _08151_ _09096_ vssd1 vssd1 vccd1 vccd1 _09226_ sky130_fd_sc_hd__o22ai_1
XFILLER_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13795_ _06057_ _06530_ _06531_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__o21ba_1
X_18322_ _02020_ _02021_ _09817_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__o21a_1
X_15534_ _08170_ _08178_ vssd1 vssd1 vccd1 vccd1 _08179_ sky130_fd_sc_hd__nor2_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12746_ _05492_ _05493_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__or2_2
XFILLER_203_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18253_ _01859_ _01863_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__nand2_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15465_ _08109_ _08085_ _08104_ vssd1 vssd1 vccd1 vccd1 _08110_ sky130_fd_sc_hd__or3_1
XFILLER_129_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12677_ rbzero.debug_overlay.facingX\[-8\] rbzero.wall_tracer.rayAddendX\[0\] vssd1
+ vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__nor2_1
XFILLER_129_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17204_ rbzero.wall_tracer.mapX\[7\] _05512_ _09782_ vssd1 vssd1 vccd1 vccd1 _09787_
+ sky130_fd_sc_hd__o21a_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14416_ _07147_ _07152_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18184_ _10271_ _01766_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__o21bai_1
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11628_ _04405_ _04406_ _04218_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__mux2_1
XFILLER_191_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15396_ _08039_ _08040_ vssd1 vssd1 vccd1 vccd1 _08041_ sky130_fd_sc_hd__nand2_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17135_ _07831_ vssd1 vssd1 vccd1 vccd1 _09763_ sky130_fd_sc_hd__buf_2
XFILLER_129_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14347_ _07059_ _07083_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__nand2_1
X_11559_ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__clkbuf_4
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17066_ _03953_ _09283_ _08377_ _09433_ vssd1 vssd1 vccd1 vccd1 _09706_ sky130_fd_sc_hd__or4_1
XFILLER_116_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14278_ _07013_ _07014_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__xor2_2
XFILLER_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16017_ _08659_ _08661_ vssd1 vssd1 vccd1 vccd1 _08662_ sky130_fd_sc_hd__nand2_1
XFILLER_83_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13229_ _05648_ _05792_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__nor2_1
XFILLER_100_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17968_ _01441_ _01547_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__or2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19707_ _03080_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16919_ _07602_ _09283_ _05209_ _09287_ vssd1 vssd1 vccd1 vccd1 _09560_ sky130_fd_sc_hd__or4_1
XFILLER_77_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17899_ _01592_ _01601_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__xnor2_1
XFILLER_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03307_ _03307_ vssd1 vssd1 vccd1 vccd1 clknet_0__03307_ sky130_fd_sc_hd__clkbuf_16
X_19638_ clknet_1_1__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__buf_1
XFILLER_93_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19569_ rbzero.pov.spi_counter\[6\] _03034_ _03036_ vssd1 vssd1 vccd1 vccd1 _00828_
+ sky130_fd_sc_hd__o21a_1
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21600_ net141 _01369_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21531_ net452 _01300_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21462_ net383 _01231_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20413_ rbzero.traced_texa\[-12\] rbzero.texV\[-12\] vssd1 vssd1 vccd1 vccd1 _03325_
+ sky130_fd_sc_hd__nand2_1
XFILLER_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21393_ net314 _01162_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20352__361 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__inv_2
XFILLER_107_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10930_ rbzero.tex_b1\[26\] rbzero.tex_b1\[27\] _03806_ vssd1 vssd1 vccd1 vccd1 _03812_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10861_ rbzero.tex_b1\[59\] rbzero.tex_b1\[60\] _03773_ vssd1 vssd1 vccd1 vccd1 _03776_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12600_ rbzero.debug_overlay.facingY\[-9\] rbzero.wall_tracer.rayAddendY\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__or2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _06287_ _06286_ _05988_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__o21a_1
XFILLER_12_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10792_ _03739_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__clkbuf_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _05285_ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_157_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15250_ _07595_ _07592_ vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__nand2_1
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12462_ rbzero.wall_tracer.trackDistX\[8\] vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__inv_2
XFILLER_8_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14201_ _06805_ _06678_ _06937_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__or3b_1
X_11413_ rbzero.row_render.size\[2\] gpout0.hpos\[2\] _04163_ gpout0.hpos\[0\] vssd1
+ vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__a22o_1
Xtop_ew_algofoogle_82 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_82/HI o_rgb[12] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_93 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_93/HI zeros[3] sky130_fd_sc_hd__conb_1
X_15181_ _07820_ _04462_ _07833_ _07834_ vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__o22ai_1
X_12393_ _05145_ _05143_ _04021_ _05159_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__a31o_1
XFILLER_138_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _06863_ _06868_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11344_ _04082_ _04088_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__nand2_1
XFILLER_192_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14063_ _06786_ _06794_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__xor2_1
X_18940_ _02599_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] vssd1 vssd1
+ vccd1 vccd1 _04055_ sky130_fd_sc_hd__nand2_1
XFILLER_180_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13014_ _05750_ _05702_ _05683_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__or3_1
X_18871_ rbzero.wall_tracer.trackDistY\[10\] rbzero.wall_tracer.stepDistY\[10\] vssd1
+ vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__or2_1
XFILLER_67_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17822_ _01524_ _01525_ _10131_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__or3b_1
XFILLER_95_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 rbzero.pov.spi_buffer\[31\] vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17753_ _10235_ _10253_ _01456_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__a21o_1
X_14965_ _07652_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_48_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16704_ _09220_ _09344_ vssd1 vssd1 vccd1 vccd1 _09346_ sky130_fd_sc_hd__and2_1
X_20180__206 clknet_1_0__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__inv_2
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13916_ _06644_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__xnor2_1
X_17684_ _09670_ _10099_ vssd1 vssd1 vccd1 vccd1 _10249_ sky130_fd_sc_hd__nand2_1
X_14896_ _07591_ _07604_ _07605_ _04039_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__o211a_1
XFILLER_130_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16635_ _08242_ _09129_ _08180_ vssd1 vssd1 vccd1 vccd1 _09278_ sky130_fd_sc_hd__a21oi_1
X_19423_ _02906_ rbzero.wall_tracer.rayAddendY\[2\] vssd1 vssd1 vccd1 vccd1 _02907_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _06263_ _06582_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__and2_1
XFILLER_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16566_ _09175_ _09176_ _09178_ vssd1 vssd1 vccd1 vccd1 _09209_ sky130_fd_sc_hd__o21ai_1
XFILLER_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19354_ _02840_ _02841_ _02842_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__o21ai_1
X_13778_ _06513_ _06514_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__and2b_1
XFILLER_206_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18305_ _02003_ _02004_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__and2b_1
X_15517_ _08135_ vssd1 vssd1 vccd1 vccd1 _08162_ sky130_fd_sc_hd__clkbuf_4
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12729_ _05424_ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__and2_1
X_19285_ _02797_ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__clkbuf_1
X_16497_ _08985_ vssd1 vssd1 vccd1 vccd1 _09141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18236_ _01933_ _01935_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__nand2_1
XFILLER_50_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15448_ _08028_ _08092_ vssd1 vssd1 vccd1 vccd1 _08093_ sky130_fd_sc_hd__and2_1
XFILLER_176_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18167_ _01866_ _01867_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15379_ _07913_ _07924_ _07941_ _07967_ vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__or4_1
XFILLER_50_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17118_ _09753_ _04319_ _09754_ vssd1 vssd1 vccd1 vccd1 _09755_ sky130_fd_sc_hd__and3_1
XFILLER_143_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18098_ _01670_ _01673_ _01789_ _01669_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__a211o_1
XFILLER_172_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17049_ _09683_ _09688_ vssd1 vssd1 vccd1 vccd1 _09689_ sky130_fd_sc_hd__and2_1
XFILLER_143_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20962_ clknet_leaf_7_i_clk _00731_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893_ clknet_leaf_86_i_clk _00662_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21514_ net435 _01283_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20276__292 clknet_1_1__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__inv_2
XFILLER_182_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21445_ net366 _01214_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21376_ net297 _01145_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20327_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__buf_1
XFILLER_162_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11060_ rbzero.tex_b0\[29\] rbzero.tex_b0\[28\] _03876_ vssd1 vssd1 vccd1 vccd1 _03880_
+ sky130_fd_sc_hd__mux2_1
XFILLER_118_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ rbzero.wall_tracer.stepDistY\[-10\] _07484_ _07461_ vssd1 vssd1 vccd1 vccd1
+ _07485_ sky130_fd_sc_hd__mux2_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11962_ _04735_ _04737_ _04324_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__o21bai_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _06436_ _06437_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__nand2_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ rbzero.tex_b1\[34\] rbzero.tex_b1\[35\] _03795_ vssd1 vssd1 vccd1 vccd1 _03803_
+ sky130_fd_sc_hd__mux2_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14681_ _07106_ _07415_ _07416_ _07417_ _05892_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__o311a_1
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _04272_ vssd1 vssd1 vccd1 vccd1 _04669_
+ sky130_fd_sc_hd__mux2_1
X_16420_ _09061_ _09062_ _09063_ vssd1 vssd1 vccd1 vccd1 _09065_ sky130_fd_sc_hd__a21o_1
X_13632_ _06352_ _06367_ _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__a21o_1
X_10844_ rbzero.tex_g0\[4\] rbzero.tex_g0\[3\] _03762_ vssd1 vssd1 vccd1 vccd1 _03767_
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16351_ _08249_ _08280_ vssd1 vssd1 vccd1 vccd1 _08996_ sky130_fd_sc_hd__nor2_1
X_13563_ _06291_ _06298_ _06299_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__o21a_1
XFILLER_157_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10775_ rbzero.tex_g0\[37\] rbzero.tex_g0\[36\] _03729_ vssd1 vssd1 vccd1 vccd1 _03731_
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15302_ rbzero.debug_overlay.playerX\[-5\] _07898_ rbzero.debug_overlay.playerX\[-4\]
+ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__o21ai_1
XFILLER_197_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19070_ _02667_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__clkbuf_1
X_12514_ rbzero.wall_tracer.trackDistY\[3\] _05264_ rbzero.wall_tracer.trackDistY\[2\]
+ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__o22a_1
X_16282_ _08924_ _08926_ vssd1 vssd1 vccd1 vccd1 _08927_ sky130_fd_sc_hd__nor2_1
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13494_ _06196_ _06230_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__xnor2_1
XFILLER_173_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18021_ _01722_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__inv_2
XFILLER_173_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15233_ _07870_ _07873_ _07881_ _07830_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__a31o_1
XFILLER_201_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12445_ _05201_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__clkbuf_4
XFILLER_154_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15164_ _07788_ _07797_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__nand2_1
X_12376_ net32 vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__clkbuf_4
XFILLER_5_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14115_ _06675_ _06690_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__nor2_1
XFILLER_5_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11327_ _04101_ _04105_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__o21ba_1
XFILLER_180_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19972_ rbzero.pov.ready_buffer\[23\] _03240_ _03243_ rbzero.debug_overlay.facingY\[-8\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__o221a_1
X_15095_ _07703_ _07753_ _07754_ _07706_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__a31o_1
XFILLER_119_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18923_ _02588_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__clkbuf_1
X_14046_ _06781_ _06782_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__or2b_1
X_11258_ _04035_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__buf_4
XFILLER_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18854_ _02529_ _02016_ rbzero.wall_tracer.trackDistY\[7\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00620_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11189_ _03977_ _03936_ _03919_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__and3b_1
X_17805_ _09276_ _09674_ _10245_ _01508_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__o31a_1
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18785_ _02468_ _05531_ _02469_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__or3b_1
X_15997_ _07598_ _07951_ _05207_ _07927_ vssd1 vssd1 vccd1 vccd1 _08642_ sky130_fd_sc_hd__or4b_2
XFILLER_94_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17736_ _10285_ _10287_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__nor2_1
XFILLER_35_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14948_ _04035_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__clkbuf_4
XFILLER_36_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17667_ _10199_ _10231_ vssd1 vssd1 vccd1 vccd1 _10232_ sky130_fd_sc_hd__xnor2_1
X_14879_ _05278_ vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__buf_4
XFILLER_165_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19406_ _04035_ _02882_ _02891_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__a21o_1
X_16618_ _09259_ _09260_ vssd1 vssd1 vccd1 vccd1 _09261_ sky130_fd_sc_hd__nor2_1
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17598_ _10039_ _10163_ vssd1 vssd1 vccd1 vccd1 _10164_ sky130_fd_sc_hd__xnor2_1
XFILLER_206_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16549_ _09089_ _09192_ vssd1 vssd1 vccd1 vccd1 _09193_ sky130_fd_sc_hd__xnor2_2
X_19337_ rbzero.debug_overlay.vplaneY\[-7\] rbzero.wall_tracer.rayAddendY\[-7\] vssd1
+ vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__nor2_1
XFILLER_204_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19268_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_floor\[4\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__mux2_1
XFILLER_148_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18219_ _01854_ _01819_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__or2b_1
X_19199_ rbzero.spi_registers.new_sky\[3\] rbzero.color_sky\[3\] _02740_ vssd1 vssd1
+ vccd1 vccd1 _02746_ sky130_fd_sc_hd__mux2_1
XFILLER_141_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21230_ clknet_leaf_18_i_clk _00999_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21161_ clknet_leaf_84_i_clk _00930_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21092_ net182 _00861_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20043_ _04887_ _04886_ _03278_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__and3_1
XFILLER_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ clknet_leaf_5_i_clk _00714_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20876_ clknet_leaf_97_i_clk _00645_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10560_ _03617_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _03581_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12230_ gpout2.clk_div\[1\] _04981_ _04999_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21428_ net349 _01197_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12161_ gpout0.hpos\[0\] _04163_ _04910_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__mux2_1
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_31_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_21359_ net280 _01128_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11112_ rbzero.tex_b0\[4\] rbzero.tex_b0\[3\] _03898_ vssd1 vssd1 vccd1 vccd1 _03907_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12092_ _04021_ _04855_ _04853_ net42 vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__a22o_1
XFILLER_104_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15920_ _08564_ _08503_ vssd1 vssd1 vccd1 vccd1 _08565_ sky130_fd_sc_hd__xor2_1
X_11043_ rbzero.tex_b0\[37\] rbzero.tex_b0\[36\] _03865_ vssd1 vssd1 vccd1 vccd1 _03871_
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_15851_ _08495_ _08141_ vssd1 vssd1 vccd1 vccd1 _08496_ sky130_fd_sc_hd__xnor2_1
XFILLER_7_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _07473_ _07492_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__nand2_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18570_ _02265_ _02266_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__xnor2_1
X_15782_ _08425_ vssd1 vssd1 vccd1 vccd1 _08427_ sky130_fd_sc_hd__clkbuf_4
XFILLER_58_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _05702_ _05729_ _05730_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__nor3_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17521_ _10085_ _10086_ vssd1 vssd1 vccd1 vccd1 _10087_ sky130_fd_sc_hd__nand2_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ _07467_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__clkbuf_4
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ rbzero.tex_b0\[46\] _04337_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__and2_1
XFILLER_91_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17452_ _09918_ _10018_ vssd1 vssd1 vccd1 vccd1 _10019_ sky130_fd_sc_hd__xnor2_4
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _05893_ _07041_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__and2_1
X_11876_ rbzero.tex_g1\[27\] rbzero.tex_g1\[26\] _04271_ vssd1 vssd1 vccd1 vccd1 _04653_
+ sky130_fd_sc_hd__mux2_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16403_ _08165_ _08432_ vssd1 vssd1 vccd1 vccd1 _09048_ sky130_fd_sc_hd__and2_2
X_13615_ _06338_ _06343_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__xnor2_1
X_17383_ _09947_ _09949_ vssd1 vssd1 vccd1 vccd1 _09950_ sky130_fd_sc_hd__xor2_1
XFILLER_60_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10827_ rbzero.tex_g0\[12\] rbzero.tex_g0\[11\] _03751_ vssd1 vssd1 vccd1 vccd1 _03758_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14595_ _07216_ _07331_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__and2_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16334_ _08977_ _08978_ vssd1 vssd1 vccd1 vccd1 _08979_ sky130_fd_sc_hd__xnor2_2
X_19122_ net42 rbzero.spi_registers.mosi_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02696_ sky130_fd_sc_hd__mux2_1
X_20292__307 clknet_1_1__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__inv_2
X_13546_ _05824_ _06080_ _06282_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__or3_2
X_10758_ rbzero.tex_g0\[45\] rbzero.tex_g0\[44\] _03718_ vssd1 vssd1 vccd1 vccd1 _03722_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19053_ _02658_ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__clkbuf_1
X_16265_ _08901_ _08908_ _08909_ vssd1 vssd1 vccd1 vccd1 _08910_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13477_ _06041_ _06067_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__or2_1
X_10689_ _03685_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18004_ _08445_ _09353_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__nand2_1
X_15216_ _07863_ _07867_ _00013_ rbzero.wall_tracer.rayAddendX\[8\] vssd1 vssd1 vccd1
+ vccd1 _00504_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12428_ net71 rbzero.wall_tracer.state\[12\] _05190_ vssd1 vssd1 vccd1 vccd1 _05191_
+ sky130_fd_sc_hd__and3_1
XFILLER_173_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16196_ _08831_ _08837_ _08839_ vssd1 vssd1 vccd1 vccd1 _08841_ sky130_fd_sc_hd__and3_1
XFILLER_142_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15147_ _07730_ rbzero.debug_overlay.vplaneX\[-5\] _07800_ _07801_ vssd1 vssd1 vccd1
+ vccd1 _07803_ sky130_fd_sc_hd__nor4_1
XFILLER_99_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12359_ gpout4.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__clkinv_2
XFILLER_5_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15078_ rbzero.debug_overlay.vplaneX\[-6\] _07735_ _07738_ vssd1 vssd1 vccd1 vccd1
+ _07739_ sky130_fd_sc_hd__o21ai_1
X_19955_ _02721_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__buf_2
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18906_ rbzero.spi_registers.spi_counter\[0\] _02558_ vssd1 vssd1 vccd1 vccd1 _02576_
+ sky130_fd_sc_hd__nand2_1
X_14029_ _06762_ _06764_ _06765_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__nand3_1
XFILLER_101_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19886_ _03192_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__clkbuf_4
XFILLER_171_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18837_ _02513_ _02514_ _01792_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__o21ai_1
XFILLER_56_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18768_ _09812_ _02454_ _09877_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__o21ai_1
X_17719_ _10281_ _10283_ vssd1 vssd1 vccd1 vccd1 _10284_ sky130_fd_sc_hd__xor2_1
XFILLER_64_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18699_ _02390_ _02394_ rbzero.wall_tracer.trackDistX\[11\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00600_ sky130_fd_sc_hd__o2bb2a_1
X_20730_ clknet_leaf_84_i_clk _00499_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20661_ clknet_leaf_63_i_clk _00445_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_91_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20592_ _02829_ _02831_ _02830_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__a21bo_1
XFILLER_177_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21213_ clknet_leaf_26_i_clk _00982_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21144_ clknet_leaf_97_i_clk _00913_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21075_ net165 _00844_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_150_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20026_ _03259_ _03268_ _03269_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__a21oi_1
XFILLER_150_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11730_ rbzero.debug_overlay.playerX\[-6\] _04475_ _04454_ rbzero.debug_overlay.playerX\[-5\]
+ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__a22o_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20928_ clknet_leaf_26_i_clk _00697_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _04418_ _04430_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__and2_1
X_20859_ clknet_leaf_2_i_clk _00628_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ _06068_ _06064_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__xor2_1
X_10612_ _03644_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__clkbuf_1
X_14380_ _06176_ _07116_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__and2_1
X_11592_ _04119_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__buf_4
X_13331_ _06065_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__nor2_1
X_10543_ _03608_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16050_ _08692_ _08694_ vssd1 vssd1 vccd1 vccd1 _08695_ sky130_fd_sc_hd__nor2_2
X_13262_ _05977_ _05987_ _05997_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__and3_1
XFILLER_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10474_ _03572_ vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15001_ rbzero.wall_tracer.stepDistX\[7\] _07575_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07671_ sky130_fd_sc_hd__mux2_1
X_12213_ _04977_ net16 _04979_ _04982_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__a31o_1
XFILLER_108_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ _05901_ _05891_ _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__a21oi_1
XFILLER_155_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20135__166 clknet_1_0__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__inv_2
XFILLER_123_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12144_ _04910_ _04325_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__nor2_1
XFILLER_150_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19740_ rbzero.pov.spi_buffer\[44\] rbzero.pov.spi_buffer\[45\] _03092_ vssd1 vssd1
+ vccd1 vccd1 _03098_ sky130_fd_sc_hd__mux2_1
X_12075_ _04840_ _04738_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__nor2_1
X_16952_ _09454_ _09591_ vssd1 vssd1 vccd1 vccd1 _09593_ sky130_fd_sc_hd__nor2_1
XFILLER_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15903_ _08470_ _08546_ vssd1 vssd1 vccd1 vccd1 _08548_ sky130_fd_sc_hd__and2_1
X_11026_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _03854_ vssd1 vssd1 vccd1 vccd1 _03862_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19671_ rbzero.pov.spi_buffer\[11\] rbzero.pov.spi_buffer\[12\] _03059_ vssd1 vssd1
+ vccd1 vccd1 _03062_ sky130_fd_sc_hd__mux2_1
X_16883_ _09521_ _09523_ vssd1 vssd1 vccd1 vccd1 _09524_ sky130_fd_sc_hd__nand2_1
X_18622_ _02317_ _02318_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__nand2_1
XFILLER_92_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _08477_ _08472_ vssd1 vssd1 vccd1 vccd1 _08479_ sky130_fd_sc_hd__xor2_2
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18553_ _02235_ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__xnor2_1
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _08372_ _08399_ vssd1 vssd1 vccd1 vccd1 _08410_ sky130_fd_sc_hd__nor2_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12977_ _05567_ _05599_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__nor2_2
XFILLER_166_1120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17504_ _09391_ _08427_ _09941_ _09942_ vssd1 vssd1 vccd1 vccd1 _10070_ sky130_fd_sc_hd__o31ai_2
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11928_ rbzero.tex_b0\[57\] _04327_ _04328_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__and3_1
XFILLER_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14716_ _07104_ _07450_ _07451_ _07452_ _05742_ _07375_ vssd1 vssd1 vccd1 vccd1 _07453_
+ sky130_fd_sc_hd__mux4_2
X_18484_ _02171_ _02181_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__nand2_1
X_15696_ _08338_ _08339_ vssd1 vssd1 vccd1 vccd1 _08341_ sky130_fd_sc_hd__nand2_1
XFILLER_205_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20300__314 clknet_1_1__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__inv_2
XFILLER_162_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17435_ _10000_ _10001_ vssd1 vssd1 vccd1 vccd1 _10002_ sky130_fd_sc_hd__xnor2_2
XFILLER_33_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14647_ _05893_ _07101_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__nor2_1
X_11859_ _04379_ _04633_ _04634_ _04635_ _04229_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__o221a_1
XFILLER_127_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_18 _09162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _09931_ _09932_ vssd1 vssd1 vccd1 vccd1 _09933_ sky130_fd_sc_hd__or2_1
X_14578_ _07311_ _07313_ _07314_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__a21o_1
XFILLER_119_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19105_ rbzero.spi_registers.spi_buffer\[8\] rbzero.spi_registers.spi_buffer\[7\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__mux2_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16317_ _07924_ _08276_ vssd1 vssd1 vccd1 vccd1 _08962_ sky130_fd_sc_hd__nor2_1
XFILLER_118_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13529_ _06255_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__xnor2_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17297_ _09807_ _09194_ vssd1 vssd1 vccd1 vccd1 _09869_ sky130_fd_sc_hd__or2_1
XFILLER_174_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16248_ _08872_ _08128_ _08868_ vssd1 vssd1 vccd1 vccd1 _08893_ sky130_fd_sc_hd__or3_1
X_19036_ rbzero.pov.spi_buffer\[49\] rbzero.pov.ready_buffer\[49\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02650_ sky130_fd_sc_hd__mux2_1
XFILLER_174_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16179_ _08519_ _08823_ _08329_ _08377_ vssd1 vssd1 vccd1 vccd1 _08824_ sky130_fd_sc_hd__o22ai_1
XFILLER_115_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19938_ _03920_ _03227_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__and2_1
XFILLER_29_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19869_ rbzero.debug_overlay.playerX\[2\] _03155_ _03179_ _03157_ vssd1 vssd1 vccd1
+ vccd1 _00985_ sky130_fd_sc_hd__o211a_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20713_ clknet_leaf_62_i_clk _00004_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20644_ clknet_leaf_59_i_clk _00428_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
X_20575_ gpout1.clk_div\[0\] gpout1.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__nand2_1
XFILLER_178_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21127_ clknet_leaf_94_i_clk _00896_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21058_ clknet_leaf_0_i_clk _00827_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_143_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12900_ _05628_ _05626_ _05633_ _05631_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__a211o_1
X_20009_ _03256_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_101_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13880_ _06592_ _06567_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__and2b_1
XFILLER_47_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ rbzero.wall_tracer.visualWallDist\[8\] _04031_ vssd1 vssd1 vccd1 vccd1 _05568_
+ sky130_fd_sc_hd__nor2_1
XFILLER_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15550_ _07893_ _05369_ vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__nor2_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ rbzero.debug_overlay.playerX\[2\] _05508_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05509_ sky130_fd_sc_hd__mux2_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14501_ _06002_ _07072_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__nand2_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11713_ rbzero.debug_overlay.facingX\[0\] _04459_ _04460_ rbzero.debug_overlay.facingX\[-2\]
+ _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__a221o_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _08034_ _08046_ _08124_ _08125_ vssd1 vssd1 vccd1 vccd1 _08126_ sky130_fd_sc_hd__or4_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _05436_ _05440_ _05434_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__o21a_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _07141_ _07140_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__and2b_1
X_17220_ rbzero.wall_tracer.mapX\[10\] _05525_ _09799_ vssd1 vssd1 vccd1 vccd1 _09800_
+ sky130_fd_sc_hd__a21bo_1
X_11644_ _04415_ _04417_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__and2b_1
XFILLER_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17151_ rbzero.row_render.texu\[1\] _09766_ _07728_ rbzero.wall_tracer.texu\[1\]
+ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__a22o_1
XFILLER_122_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14363_ _07043_ _07098_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__nor2_1
X_11575_ _04306_ _04346_ _04353_ _04241_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__a211o_1
Xinput16 i_gpout2_sel[2] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__buf_8
XFILLER_196_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput27 i_gpout4_sel[1] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16102_ _07601_ _08227_ vssd1 vssd1 vccd1 vccd1 _08747_ sky130_fd_sc_hd__nand2_2
XFILLER_122_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput38 i_mode[0] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_8
X_13314_ _06021_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__xnor2_1
Xinput49 i_tex_in[3] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_4
X_10526_ _03599_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__clkbuf_1
X_17082_ _09680_ _09721_ vssd1 vssd1 vccd1 vccd1 _09722_ sky130_fd_sc_hd__xnor2_2
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14294_ _06735_ _07030_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__xnor2_2
XFILLER_196_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16033_ _08676_ _08677_ vssd1 vssd1 vccd1 vccd1 _08678_ sky130_fd_sc_hd__and2_1
XFILLER_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ _05981_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__clkbuf_4
X_10457_ _03563_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ _05778_ _05829_ _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__a21o_1
X_10388_ rbzero.tex_r1\[25\] rbzero.tex_r1\[26\] _03516_ vssd1 vssd1 vccd1 vccd1 _03525_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12127_ _04851_ _04896_ _04898_ _04865_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__a22o_2
XFILLER_124_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17984_ _01445_ _01447_ _01571_ _01569_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__a31o_1
X_19723_ rbzero.pov.spi_buffer\[36\] rbzero.pov.spi_buffer\[37\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03089_ sky130_fd_sc_hd__mux2_1
X_12058_ _04812_ _04817_ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__or3b_1
X_16935_ _09439_ _09440_ vssd1 vssd1 vccd1 vccd1 _09576_ sky130_fd_sc_hd__nor2_1
XFILLER_133_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11009_ rbzero.tex_b0\[53\] rbzero.tex_b0\[52\] _03843_ vssd1 vssd1 vccd1 vccd1 _03853_
+ sky130_fd_sc_hd__mux2_1
XFILLER_133_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19654_ rbzero.pov.spi_buffer\[3\] rbzero.pov.spi_buffer\[4\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03053_ sky130_fd_sc_hd__mux2_1
XFILLER_65_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16866_ _09499_ _09506_ vssd1 vssd1 vccd1 vccd1 _09507_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18605_ _02204_ _02214_ _02202_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a21oi_1
XFILLER_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15817_ _08441_ _08459_ vssd1 vssd1 vccd1 vccd1 _08462_ sky130_fd_sc_hd__nor2_1
XFILLER_93_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16797_ _09425_ _09438_ vssd1 vssd1 vccd1 vccd1 _09439_ sky130_fd_sc_hd__xnor2_2
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18536_ _02232_ _02233_ _09817_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__o21a_1
X_15748_ _07996_ _08194_ _08386_ _08385_ vssd1 vssd1 vccd1 vccd1 _08393_ sky130_fd_sc_hd__o31a_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18467_ _02054_ _02035_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__or2b_1
X_15679_ _08317_ _08323_ vssd1 vssd1 vccd1 vccd1 _08324_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17418_ _09979_ _09984_ vssd1 vssd1 vccd1 vccd1 _09985_ sky130_fd_sc_hd__xor2_2
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18398_ _02093_ _02095_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__nand2_1
XFILLER_202_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17349_ _09654_ _09909_ _09914_ vssd1 vssd1 vccd1 vccd1 _09916_ sky130_fd_sc_hd__and3_1
XFILLER_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20360_ clknet_1_0__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__buf_1
XFILLER_162_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19019_ rbzero.pov.spi_buffer\[41\] rbzero.pov.ready_buffer\[41\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02641_ sky130_fd_sc_hd__mux2_1
X_20118__150 clknet_1_0__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__inv_2
XFILLER_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19587__43 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__inv_2
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03312_ clknet_0__03312_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03312_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20627_ clknet_leaf_17_i_clk _00411_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_col\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_153_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11360_ _04116_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__clkinv_4
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20558_ _09763_ _09859_ rbzero.traced_texVinit\[2\] _09762_ vssd1 vssd1 vccd1 vccd1
+ _01410_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_180_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10311_ rbzero.tex_r1\[62\] rbzero.tex_r1\[63\] _03483_ vssd1 vssd1 vccd1 vccd1 _03485_
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11291_ rbzero.texV\[5\] _04070_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__xor2_1
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20489_ _03272_ _03386_ _03388_ _03250_ rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1
+ _01396_ sky130_fd_sc_hd__a32o_1
XFILLER_152_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13030_ _05725_ _05764_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a21bo_1
XFILLER_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14981_ rbzero.wall_tracer.stepDistX\[-3\] _07545_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07661_ sky130_fd_sc_hd__mux2_1
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16720_ _09352_ _09361_ vssd1 vssd1 vccd1 vccd1 _09362_ sky130_fd_sc_hd__xnor2_1
X_13932_ _06659_ _06664_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20247__267 clknet_1_0__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__inv_2
XFILLER_75_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16651_ _05211_ _09138_ vssd1 vssd1 vccd1 vccd1 _09294_ sky130_fd_sc_hd__or2_2
X_13863_ _06335_ _06560_ _06562_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__and3_1
XFILLER_207_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15602_ _08242_ _08239_ _08245_ _08246_ vssd1 vssd1 vccd1 vccd1 _08247_ sky130_fd_sc_hd__o31a_2
X_12814_ _05533_ _05551_ _05553_ _05284_ rbzero.wall_tracer.mapY\[9\] vssd1 vssd1
+ vccd1 vccd1 _00416_ sky130_fd_sc_hd__a32o_1
X_19370_ rbzero.wall_tracer.rayAddendY\[-3\] _02858_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _02859_ sky130_fd_sc_hd__mux2_1
X_16582_ _08821_ _08823_ _08419_ vssd1 vssd1 vccd1 vccd1 _09225_ sky130_fd_sc_hd__or3_1
X_13794_ _06511_ _06512_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__nand2_1
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18321_ _02017_ _02018_ _02019_ _05531_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__a31o_1
X_15533_ _08177_ vssd1 vssd1 vccd1 vccd1 _08178_ sky130_fd_sc_hd__clkbuf_4
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _05446_ _05447_ _05451_ _05449_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__o211a_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18252_ _01841_ _01842_ _01844_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__a21bo_1
X_15464_ _08074_ vssd1 vssd1 vccd1 vccd1 _08109_ sky130_fd_sc_hd__clkbuf_4
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__nand2_2
XFILLER_163_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14415_ _07132_ _07151_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__xnor2_1
X_17203_ rbzero.wall_tracer.mapX\[7\] _09781_ _09779_ _09786_ vssd1 vssd1 vccd1 vccd1
+ _00572_ sky130_fd_sc_hd__a22o_1
X_11627_ rbzero.tex_r1\[37\] rbzero.tex_r1\[36\] _04250_ vssd1 vssd1 vccd1 vccd1 _04406_
+ sky130_fd_sc_hd__mux2_1
X_18183_ _01646_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15395_ _05197_ rbzero.wall_tracer.stepDistX\[-9\] vssd1 vssd1 vccd1 vccd1 _08040_
+ sky130_fd_sc_hd__or2_1
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14346_ _07080_ _07082_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__xor2_1
X_17134_ rbzero.row_render.side _09762_ _07728_ _07895_ vssd1 vssd1 vccd1 vccd1 _00527_
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11558_ _04336_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__buf_6
XFILLER_183_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10509_ _03590_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__clkbuf_1
X_17065_ _07602_ _09283_ _05210_ _09433_ vssd1 vssd1 vccd1 vccd1 _09705_ sky130_fd_sc_hd__or4_1
XFILLER_128_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14277_ _06689_ _06668_ _06750_ _06748_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__o31a_1
XFILLER_109_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11489_ _04244_ _04256_ _04268_ _04116_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a31o_1
XFILLER_48_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16016_ _08574_ _08660_ vssd1 vssd1 vccd1 vccd1 _08661_ sky130_fd_sc_hd__and2_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ _05697_ _05792_ _05778_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__a21o_1
XFILLER_83_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _05802_ _05815_ _05884_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__mux2_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _10183_ _09906_ _10294_ _01550_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__or4bb_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19706_ rbzero.pov.spi_buffer\[28\] rbzero.pov.spi_buffer\[29\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03080_ sky130_fd_sc_hd__mux2_1
XFILLER_78_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16918_ _09553_ _09558_ vssd1 vssd1 vccd1 vccd1 _09559_ sky130_fd_sc_hd__xnor2_2
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17898_ _01599_ _01600_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__and2b_1
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03306_ _03306_ vssd1 vssd1 vccd1 vccd1 clknet_0__03306_ sky130_fd_sc_hd__clkbuf_16
X_19637_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__buf_1
X_16849_ _08823_ _09164_ _09354_ vssd1 vssd1 vccd1 vccd1 _09490_ sky130_fd_sc_hd__or3_1
XFILLER_66_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19568_ rbzero.pov.spi_counter\[6\] _03034_ _03026_ vssd1 vssd1 vccd1 vccd1 _03036_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18519_ _02105_ _02115_ _02216_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__a21oi_1
XFILLER_181_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19499_ _02952_ _02975_ _02976_ _02977_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__nand4_1
XFILLER_179_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21530_ net451 _01299_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21461_ net382 _01230_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[40\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_opt_9_0_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_9_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20412_ _03324_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21392_ net313 _01161_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_88_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _03775_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_186_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10791_ rbzero.tex_g0\[29\] rbzero.tex_g0\[28\] _03729_ vssd1 vssd1 vccd1 vccd1 _03739_
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _05205_ rbzero.map_rom.d6 _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__mux2_1
XFILLER_9_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _05214_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.trackDistY\[9\]
+ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_200_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21659_ clknet_leaf_80_i_clk _01428_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14200_ _06926_ _06935_ _06936_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__a21oi_1
X_11412_ rbzero.row_render.size\[0\] gpout0.hpos\[0\] _04163_ vssd1 vssd1 vccd1 vccd1
+ _04192_ sky130_fd_sc_hd__a21o_1
Xtop_ew_algofoogle_72 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_72/HI o_rgb[0] sky130_fd_sc_hd__conb_1
X_15180_ _07785_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 _07834_
+ sky130_fd_sc_hd__and2_1
X_12392_ net43 _05142_ _05144_ net42 _05158_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__a221o_1
Xtop_ew_algofoogle_83 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_83/HI o_rgb[13] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_94 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_94/HI zeros[4] sky130_fd_sc_hd__conb_1
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14131_ _06828_ _06864_ _06865_ _06867_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_4_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11343_ _04093_ _04114_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__or3_4
XFILLER_165_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14062_ _06722_ _06720_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__xnor2_1
X_11274_ rbzero.traced_texVinit\[8\] rbzero.spi_registers.vshift\[5\] vssd1 vssd1
+ vccd1 vccd1 _04054_ sky130_fd_sc_hd__or2_1
XFILLER_180_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13013_ _05601_ _05638_ _05649_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__or3_1
X_18870_ _02543_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17821_ _08263_ _08266_ _10134_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__and3_1
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5 rbzero.pov.ready_buffer\[29\] vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17752_ _10236_ _10252_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__nor2_1
XFILLER_43_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14964_ rbzero.wall_tracer.stepDistX\[-11\] _07465_ _07650_ vssd1 vssd1 vccd1 vccd1
+ _07652_ sky130_fd_sc_hd__mux2_1
X_16703_ _09220_ _09344_ vssd1 vssd1 vccd1 vccd1 _09345_ sky130_fd_sc_hd__nor2_1
XFILLER_48_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13915_ _06645_ _06651_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__xnor2_1
X_17683_ _09674_ vssd1 vssd1 vccd1 vccd1 _10248_ sky130_fd_sc_hd__clkbuf_4
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14895_ rbzero.wall_tracer.visualWallDist\[-9\] _07595_ vssd1 vssd1 vccd1 vccd1 _07605_
+ sky130_fd_sc_hd__or2_1
X_19422_ _02905_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__buf_4
X_16634_ _09117_ _09276_ vssd1 vssd1 vccd1 vccd1 _09277_ sky130_fd_sc_hd__nor2_1
XFILLER_35_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13846_ _06263_ _06582_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__nor2_1
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19353_ _02840_ _02841_ _02842_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__or3_1
X_16565_ _09188_ _09191_ vssd1 vssd1 vccd1 vccd1 _09208_ sky130_fd_sc_hd__nor2_1
X_13777_ _06477_ _06479_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__xor2_1
X_10989_ _03842_ vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18304_ _02001_ _02002_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__nand2_1
XFILLER_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15516_ _08159_ _08160_ _08152_ vssd1 vssd1 vccd1 vccd1 _08161_ sky130_fd_sc_hd__nor3_1
X_19581__38 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__inv_2
X_12728_ rbzero.debug_overlay.facingX\[-9\] rbzero.wall_tracer.rayAddendX\[-1\] vssd1
+ vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__or2_1
X_19284_ rbzero.spi_registers.spi_buffer\[4\] rbzero.spi_registers.new_leak\[4\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__mux2_1
X_16496_ _09135_ _09139_ vssd1 vssd1 vccd1 vccd1 _09140_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18235_ _01462_ _09480_ _01934_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__or3_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15447_ rbzero.debug_overlay.playerX\[-2\] _08027_ rbzero.debug_overlay.playerX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__o21ai_1
X_12659_ _05408_ rbzero.wall_tracer.mapY\[5\] _05283_ vssd1 vssd1 vccd1 vccd1 _05409_
+ sky130_fd_sc_hd__mux2_1
XFILLER_157_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18166_ _09434_ _09988_ _08802_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15378_ _07958_ _08022_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__nor2_1
XFILLER_116_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ _04814_ _03474_ _04317_ vssd1 vssd1 vccd1 vccd1 _09754_ sky130_fd_sc_hd__a21o_1
X_14329_ _07062_ _07065_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18097_ _01792_ _01798_ rbzero.wall_tracer.trackDistX\[5\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00594_ sky130_fd_sc_hd__o2bb2a_1
X_17048_ _09684_ _09687_ vssd1 vssd1 vccd1 vccd1 _09688_ sky130_fd_sc_hd__xor2_1
XFILLER_143_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18999_ _02630_ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_98_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20961_ clknet_leaf_7_i_clk _00730_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20892_ clknet_leaf_87_i_clk _00661_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21513_ net434 _01282_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21444_ net365 _01213_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21375_ net296 _01144_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ _04206_ _04736_ _04314_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__a21o_1
XFILLER_29_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _06428_ _06435_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__nand2_1
XFILLER_72_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10912_ _03802_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__clkbuf_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14680_ _07378_ _07413_ _06239_ _05779_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__a211o_1
XFILLER_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11892_ rbzero.tex_b0\[15\] _04327_ _04328_ _04329_ vssd1 vssd1 vccd1 vccd1 _04668_
+ sky130_fd_sc_hd__a31o_1
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13631_ _06366_ _06354_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__and2b_1
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10843_ _03766_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16350_ _08970_ _08994_ vssd1 vssd1 vccd1 vccd1 _08995_ sky130_fd_sc_hd__xnor2_4
XFILLER_125_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13562_ _06289_ _06290_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__nand2_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10774_ _03730_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__clkbuf_1
X_20359__368 clknet_1_1__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__inv_2
XFILLER_13_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15301_ rbzero.debug_overlay.playerX\[-4\] rbzero.debug_overlay.playerX\[-5\] _07898_
+ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__or3_1
X_12513_ rbzero.wall_tracer.trackDistX\[2\] vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__inv_2
XFILLER_158_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16281_ _08915_ _08925_ _08921_ vssd1 vssd1 vccd1 vccd1 _08926_ sky130_fd_sc_hd__o21a_1
XFILLER_73_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13493_ _06227_ _06229_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__xor2_1
XFILLER_200_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18020_ _01720_ _01721_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15232_ _07870_ _07873_ _07881_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__a21oi_1
X_12444_ _05200_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__buf_2
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ _07816_ _07817_ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__nand2_1
X_12375_ _05141_ net32 vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__and2_1
XFILLER_153_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14114_ _06848_ _06850_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11326_ _04103_ _04104_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__nor2_1
X_15094_ _07738_ _07752_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__nand2_1
XFILLER_4_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19971_ rbzero.pov.ready_buffer\[22\] _03240_ _03243_ rbzero.debug_overlay.facingY\[-9\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__o221a_1
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18922_ _02574_ _02586_ _02587_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__and3_1
XFILLER_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14045_ _06774_ _06775_ _06780_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__a21o_1
X_11257_ _04037_ rbzero.wall_tracer.state\[14\] vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__and2b_1
XFILLER_45_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18853_ _02527_ _02528_ _02406_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__o21a_1
XFILLER_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11188_ rbzero.map_rom.f3 rbzero.map_rom.f2 rbzero.map_rom.i_col\[4\] vssd1 vssd1
+ vccd1 vccd1 _03977_ sky130_fd_sc_hd__or3_1
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17804_ _10099_ _10244_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__nand2_1
XFILLER_121_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18784_ _02465_ _02466_ _02467_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__or3_1
XFILLER_95_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15996_ _08593_ _08595_ vssd1 vssd1 vccd1 vccd1 _08641_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17735_ _05268_ _09781_ _01439_ vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__a21oi_1
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14947_ rbzero.wall_tracer.visualWallDist\[7\] _07594_ vssd1 vssd1 vccd1 vccd1 _07641_
+ sky130_fd_sc_hd__or2_1
XFILLER_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17666_ _10214_ _10230_ vssd1 vssd1 vccd1 vccd1 _10231_ sky130_fd_sc_hd__xor2_1
XFILLER_169_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14878_ _04019_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__clkbuf_4
XFILLER_91_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19405_ _03913_ _02889_ _02890_ _07695_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__a31o_1
XFILLER_165_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16617_ _09256_ _09258_ vssd1 vssd1 vccd1 vccd1 _09260_ sky130_fd_sc_hd__and2_1
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13829_ _06271_ _06269_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__or2b_1
X_17597_ _10160_ _10162_ vssd1 vssd1 vccd1 vccd1 _10163_ sky130_fd_sc_hd__xor2_1
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19336_ rbzero.debug_overlay.vplaneY\[-6\] rbzero.wall_tracer.rayAddendY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__or2_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16548_ _09188_ _09191_ vssd1 vssd1 vccd1 vccd1 _09192_ sky130_fd_sc_hd__xor2_2
XFILLER_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19267_ _02787_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16479_ _09121_ _09122_ vssd1 vssd1 vccd1 vccd1 _09123_ sky130_fd_sc_hd__xnor2_1
X_18218_ _01821_ _01853_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__or2_1
XFILLER_164_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19198_ rbzero.color_sky\[2\] _02740_ _02745_ vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__a21o_1
XFILLER_15_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18149_ _01848_ _01849_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__nor2_1
XFILLER_141_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21160_ clknet_leaf_85_i_clk _00929_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_176_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21091_ net181 _00860_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20042_ _04886_ _03278_ _03280_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__o21ba_1
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20388__14 clknet_1_1__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__inv_2
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20944_ clknet_leaf_9_i_clk _00713_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20875_ clknet_leaf_96_i_clk _00644_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10490_ rbzero.tex_r0\[44\] rbzero.tex_r0\[43\] _03580_ vssd1 vssd1 vccd1 vccd1 _03581_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21427_ net348 _01196_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12160_ _04918_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__inv_2
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21358_ net279 _01127_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _03906_ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12091_ net68 _04857_ _04838_ _04323_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__a22o_1
X_21289_ clknet_leaf_37_i_clk _01058_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11042_ _03870_ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _08113_ _08139_ _08140_ vssd1 vssd1 vccd1 vccd1 _08495_ sky130_fd_sc_hd__o21bai_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _00004_ _07530_ _07531_ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__a21oi_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _08135_ _08422_ _08425_ vssd1 vssd1 vccd1 vccd1 _08426_ sky130_fd_sc_hd__or3_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12993_ _05638_ _05695_ _05677_ _05681_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__or4_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ _10051_ _10052_ _10084_ vssd1 vssd1 vccd1 vccd1 _10086_ sky130_fd_sc_hd__nand3_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _05834_ _07455_ vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__and2_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ rbzero.tex_b0\[45\] rbzero.tex_b0\[44\] _04356_ vssd1 vssd1 vccd1 vccd1 _04720_
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _10015_ _10017_ vssd1 vssd1 vccd1 vccd1 _10018_ sky130_fd_sc_hd__xnor2_2
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11875_ _04648_ _04651_ _04209_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__mux2_1
X_14663_ _07388_ _07381_ _05931_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__mux2_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _09045_ _09046_ vssd1 vssd1 vccd1 vccd1 _09047_ sky130_fd_sc_hd__nand2_2
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13614_ _06305_ _06321_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__xor2_2
XFILLER_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10826_ _03757_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__clkbuf_1
X_17382_ _09639_ _09646_ _09948_ vssd1 vssd1 vccd1 vccd1 _09949_ sky130_fd_sc_hd__a21oi_2
XFILLER_38_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14594_ _07329_ _07330_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__and2b_1
XFILLER_186_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19121_ _03555_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__buf_6
XFILLER_38_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16333_ _07598_ _08230_ _08147_ _08236_ vssd1 vssd1 vccd1 vccd1 _08978_ sky130_fd_sc_hd__or4_1
X_10757_ _03721_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__clkbuf_1
X_13545_ _06065_ _06134_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__or2_1
XFILLER_41_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19052_ rbzero.pov.spi_buffer\[57\] rbzero.pov.ready_buffer\[57\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02658_ sky130_fd_sc_hd__mux2_1
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16264_ _08897_ _08906_ _08905_ vssd1 vssd1 vccd1 vccd1 _08909_ sky130_fd_sc_hd__a21o_1
XFILLER_146_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13476_ _06179_ _06181_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__and2b_1
X_10688_ rbzero.tex_g1\[13\] rbzero.tex_g1\[14\] _03680_ vssd1 vssd1 vccd1 vccd1 _03685_
+ sky130_fd_sc_hd__mux2_1
XFILLER_139_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18003_ _01703_ _01704_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__xnor2_1
X_15215_ _07865_ _07866_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__or2_1
X_12427_ _05189_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__buf_6
X_16195_ _08831_ _08837_ _08839_ vssd1 vssd1 vccd1 vccd1 _08840_ sky130_fd_sc_hd__a21oi_1
XFILLER_138_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12358_ net52 _05103_ _05125_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__a21oi_1
XFILLER_142_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15146_ _07730_ rbzero.debug_overlay.vplaneX\[-5\] _07800_ _07801_ vssd1 vssd1 vccd1
+ vccd1 _07802_ sky130_fd_sc_hd__o22a_1
XFILLER_181_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11309_ _04082_ _04088_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__nor2_1
X_19954_ rbzero.pov.ready_buffer\[35\] _03240_ _03243_ rbzero.debug_overlay.facingX\[-7\]
+ _03209_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__o221a_1
X_15077_ rbzero.debug_overlay.vplaneX\[-6\] _07708_ _07736_ _07737_ vssd1 vssd1 vccd1
+ vccd1 _07738_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12289_ net43 _05043_ _05044_ net41 net23 vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__a221o_1
XFILLER_113_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18905_ rbzero.spi_registers.spi_counter\[0\] _02558_ vssd1 vssd1 vccd1 vccd1 _02575_
+ sky130_fd_sc_hd__or2_1
X_14028_ _05982_ _06740_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__nor2_1
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20112__145 clknet_1_1__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__inv_2
X_19885_ net39 _03137_ _02708_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__o21ai_2
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18836_ _02510_ _02511_ _02512_ _04016_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a31o_1
XFILLER_45_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18767_ _02452_ _02453_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__xnor2_1
X_15979_ _07958_ _08128_ vssd1 vssd1 vccd1 vccd1 _08624_ sky130_fd_sc_hd__nor2_1
XFILLER_49_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17718_ _10088_ _10155_ _10282_ vssd1 vssd1 vccd1 vccd1 _10283_ sky130_fd_sc_hd__a21oi_1
X_18698_ _05532_ _02393_ _09817_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__o21a_1
XFILLER_64_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17649_ _10204_ _10213_ vssd1 vssd1 vccd1 vccd1 _10214_ sky130_fd_sc_hd__xor2_1
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20660_ clknet_leaf_58_i_clk _00444_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[-11\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_205_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19319_ rbzero.spi_registers.new_vshift\[2\] rbzero.spi_registers.spi_buffer\[2\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__mux2_1
XFILLER_177_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20591_ _07679_ _02830_ _03458_ _07855_ rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__a32o_1
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21212_ clknet_leaf_26_i_clk _00981_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_145_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21143_ clknet_leaf_97_i_clk _00912_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_105_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21074_ net164 _00843_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20025_ _04892_ _04992_ _04037_ _03911_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a31o_1
XFILLER_24_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20087__122 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__inv_2
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20927_ clknet_leaf_74_i_clk _00696_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _04004_ _04438_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__and2_1
XFILLER_187_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20858_ clknet_leaf_1_i_clk _00627_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ rbzero.tex_g1\[49\] rbzero.tex_g1\[50\] _03635_ vssd1 vssd1 vccd1 vccd1 _03644_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ _04225_ _04367_ _04368_ _04369_ _04208_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__o221a_1
XFILLER_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20789_ clknet_leaf_47_i_clk _00558_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13330_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__clkbuf_4
XFILLER_195_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10542_ rbzero.tex_r0\[19\] rbzero.tex_r0\[18\] _03602_ vssd1 vssd1 vccd1 vccd1 _03608_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13261_ _05977_ _05987_ _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__a21oi_1
X_10473_ rbzero.tex_r0\[52\] rbzero.tex_r0\[51\] _03569_ vssd1 vssd1 vccd1 vccd1 _03572_
+ sky130_fd_sc_hd__mux2_1
X_12212_ net42 _04963_ _04980_ _04981_ _04021_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__a32o_1
X_15000_ _07670_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_170_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13192_ _05703_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__nor2_2
XFILLER_194_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12143_ _04910_ net64 _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__a21bo_1
XFILLER_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12074_ net5 net6 vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__nand2_1
X_16951_ _09454_ _09591_ vssd1 vssd1 vccd1 vccd1 _09592_ sky130_fd_sc_hd__and2_1
XFILLER_150_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15902_ _08470_ _08546_ vssd1 vssd1 vccd1 vccd1 _08547_ sky130_fd_sc_hd__nor2_2
X_11025_ _03861_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19670_ _03061_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16882_ _08282_ _08129_ _08047_ _09522_ vssd1 vssd1 vccd1 vccd1 _09523_ sky130_fd_sc_hd__o22ai_1
X_18621_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.stepDistX\[10\] vssd1
+ vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__nand2_1
XFILLER_49_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _08472_ _08477_ vssd1 vssd1 vccd1 vccd1 _08478_ sky130_fd_sc_hd__or2b_1
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ _02141_ _02248_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__xor2_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _08402_ _08408_ vssd1 vssd1 vccd1 vccd1 _08409_ sky130_fd_sc_hd__xnor2_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _05711_ _05712_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__xor2_2
XFILLER_166_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17503_ _10067_ _10068_ vssd1 vssd1 vccd1 vccd1 _10069_ sky130_fd_sc_hd__and2_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14715_ _07419_ _07420_ _07106_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__a21o_1
X_18483_ _02179_ _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__and2_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _04701_ _04702_ _04266_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__mux2_1
X_15695_ _08338_ _08339_ vssd1 vssd1 vccd1 vccd1 _08340_ sky130_fd_sc_hd__or2_1
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _09707_ _09708_ _09706_ vssd1 vssd1 vccd1 vccd1 _10001_ sky130_fd_sc_hd__o21a_1
XFILLER_61_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14646_ _07106_ _07379_ _07380_ _07382_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__a31o_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ rbzero.tex_g1\[10\] _04291_ _04329_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__a21o_1
XFILLER_61_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17365_ _09368_ _09165_ _09628_ _09629_ vssd1 vssd1 vccd1 vccd1 _09932_ sky130_fd_sc_hd__o31a_1
XANTENNA_19 _09350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ _03748_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__clkbuf_1
X_11789_ _04565_ _04566_ _04345_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__mux2_1
X_14577_ _07295_ _07306_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__nor2_1
XFILLER_159_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19104_ _02685_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__clkbuf_1
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16316_ _08192_ _08960_ _08179_ _08190_ vssd1 vssd1 vccd1 vccd1 _08961_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_201_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13528_ _06263_ _06264_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__and2_1
X_17296_ _09864_ _09865_ _09866_ vssd1 vssd1 vccd1 vccd1 _09868_ sky130_fd_sc_hd__a21oi_1
XFILLER_174_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19035_ _02593_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__clkbuf_4
XFILLER_173_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16247_ _08889_ _08891_ vssd1 vssd1 vccd1 vccd1 _08892_ sky130_fd_sc_hd__xor2_1
XFILLER_173_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13459_ _06194_ _06195_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__nand2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16178_ _08112_ vssd1 vssd1 vccd1 vccd1 _08823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15129_ _07785_ rbzero.wall_tracer.rayAddendX\[3\] vssd1 vssd1 vccd1 vccd1 _07786_
+ sky130_fd_sc_hd__nand2_1
XFILLER_142_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_92_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_173_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19937_ _03193_ _03230_ rbzero.debug_overlay.playerY\[4\] vssd1 vssd1 vccd1 vccd1
+ _03231_ sky130_fd_sc_hd__o21a_1
XFILLER_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19868_ rbzero.pov.ready_buffer\[70\] _02823_ _03138_ _03178_ vssd1 vssd1 vccd1 vccd1
+ _03179_ sky130_fd_sc_hd__a211o_1
XFILLER_96_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18819_ _02497_ _02498_ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__nand2_1
X_19799_ _03128_ vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03299_ clknet_0__03299_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03299_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_102_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20712_ clknet_leaf_48_i_clk _00003_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20643_ clknet_leaf_55_i_clk _00427_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20574_ gpout1.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__nor2_1
XFILLER_149_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_45_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21126_ clknet_leaf_95_i_clk _00895_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21057_ clknet_leaf_99_i_clk _00826_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20008_ _02595_ _03255_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__and2_1
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12830_ _05563_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__nand2_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _05506_ _05507_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__xor2_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _07222_ _07224_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__xnor2_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11712_ rbzero.debug_overlay.facingX\[-4\] _04464_ _04465_ rbzero.debug_overlay.facingX\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__a22o_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ rbzero.debug_overlay.facingX\[-3\] rbzero.wall_tracer.rayAddendX\[5\] vssd1
+ vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__or2_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _05196_ rbzero.wall_tracer.stepDistX\[-10\] _08053_ vssd1 vssd1 vccd1 vccd1
+ _08125_ sky130_fd_sc_hd__o21bai_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _04045_ _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__nand2_4
XFILLER_39_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _07164_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__or2_1
X_20141__171 clknet_1_1__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__inv_2
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17150_ _07706_ vssd1 vssd1 vccd1 vccd1 _09766_ sky130_fd_sc_hd__buf_4
XFILLER_196_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11574_ _04349_ _04351_ _04352_ _04225_ _04253_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__o221a_1
X_14362_ _07043_ _07098_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__and2_1
XFILLER_10_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 i_gpout2_sel[3] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_8
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16101_ _08594_ _07938_ vssd1 vssd1 vccd1 vccd1 _08746_ sky130_fd_sc_hd__nor2_1
Xinput28 i_gpout4_sel[2] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_6
Xinput39 i_mode[1] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_8
X_10525_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _03591_ vssd1 vssd1 vccd1 vccd1 _03599_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13313_ _06039_ _06048_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__o21ai_1
X_17081_ _09718_ _09720_ vssd1 vssd1 vccd1 vccd1 _09721_ sky130_fd_sc_hd__xor2_4
X_14293_ _07027_ _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__xor2_2
XFILLER_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13244_ _05941_ _05980_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__and2_1
X_16032_ _07988_ _08674_ _08020_ vssd1 vssd1 vccd1 vccd1 _08677_ sky130_fd_sc_hd__or3_1
XFILLER_115_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10456_ rbzero.tex_r0\[60\] rbzero.tex_r0\[59\] _03558_ vssd1 vssd1 vccd1 vccd1 _03563_
+ sky130_fd_sc_hd__mux2_1
XFILLER_143_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13175_ _05826_ _05911_ _05755_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__a21o_1
X_10387_ _03524_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__clkbuf_1
X_12126_ _03555_ _04857_ _04897_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__a21o_2
XFILLER_111_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17983_ _01663_ _01560_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__or2b_1
XFILLER_111_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19722_ _03088_ vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__clkbuf_1
X_12057_ _03474_ _04809_ _04810_ _04818_ _04830_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a41o_1
X_16934_ _09550_ _09574_ vssd1 vssd1 vccd1 vccd1 _09575_ sky130_fd_sc_hd__xnor2_2
XFILLER_81_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11008_ _03852_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19653_ _03052_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__clkbuf_1
X_16865_ _09500_ _09505_ vssd1 vssd1 vccd1 vccd1 _09506_ sky130_fd_sc_hd__xnor2_1
XFILLER_120_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18604_ _02291_ _02300_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__xor2_1
X_15816_ _08145_ _08122_ vssd1 vssd1 vccd1 vccd1 _08461_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16796_ _09436_ _09437_ vssd1 vssd1 vccd1 vccd1 _09438_ sky130_fd_sc_hd__xnor2_2
XFILLER_203_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18535_ _02229_ _02230_ _02231_ _05531_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__a31o_1
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20224__246 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__inv_2
X_15747_ _07943_ _07968_ _07942_ vssd1 vssd1 vccd1 vccd1 _08392_ sky130_fd_sc_hd__a21bo_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12959_ _05638_ _05682_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__or2_1
XFILLER_80_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18466_ _02083_ _02097_ _02096_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a21o_1
XFILLER_178_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15678_ _08320_ _08322_ vssd1 vssd1 vccd1 vccd1 _08323_ sky130_fd_sc_hd__xnor2_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17417_ _09982_ _09983_ vssd1 vssd1 vccd1 vccd1 _09984_ sky130_fd_sc_hd__xnor2_2
XFILLER_61_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14629_ _05793_ _07365_ vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__nand2_1
X_18397_ _02093_ _02095_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__nor2_1
XFILLER_105_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17348_ _09654_ _09909_ _09914_ vssd1 vssd1 vccd1 vccd1 _09915_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17279_ rbzero.wall_tracer.trackDistX\[-7\] _09852_ _05413_ vssd1 vssd1 vccd1 vccd1
+ _09853_ sky130_fd_sc_hd__mux2_1
XFILLER_147_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19018_ _02640_ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_175_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20270__288 clknet_1_1__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__inv_2
XFILLER_138_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_opt_5_0_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_5_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20199__223 clknet_1_0__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__inv_2
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03311_ clknet_0__03311_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03311_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20626_ clknet_leaf_16_i_clk _00410_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f1 sky130_fd_sc_hd__dfxtp_1
XFILLER_178_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20557_ rbzero.traced_texVinit\[1\] _03443_ _09771_ _09076_ vssd1 vssd1 vccd1 vccd1
+ _01409_ sky130_fd_sc_hd__a22o_1
XFILLER_193_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10310_ _03484_ vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11290_ _04067_ _04066_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__nand2_1
XFILLER_192_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20488_ _03387_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__inv_2
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21109_ net199 _00878_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[49\] sky130_fd_sc_hd__dfxtp_1
X_14980_ _05201_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__buf_4
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13931_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__clkbuf_4
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16650_ _08239_ _09292_ _09289_ _09290_ vssd1 vssd1 vccd1 vccd1 _09293_ sky130_fd_sc_hd__a2bb2o_1
X_13862_ _06277_ _06563_ _06597_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__or3b_1
XFILLER_35_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15601_ _08243_ _08244_ vssd1 vssd1 vccd1 vccd1 _08246_ sky130_fd_sc_hd__or2_1
XFILLER_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12813_ _05548_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__or2b_1
X_16581_ _09092_ _09095_ vssd1 vssd1 vccd1 vccd1 _09224_ sky130_fd_sc_hd__nand2_1
X_13793_ _05855_ _06061_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__nand2_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18320_ _02017_ _02018_ _02019_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__a21oi_1
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15532_ _08147_ rbzero.wall_tracer.stepDistX\[1\] _08175_ _08176_ vssd1 vssd1 vccd1
+ vccd1 _08177_ sky130_fd_sc_hd__a22oi_4
XFILLER_16_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[11\] vssd1
+ vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__and2_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18251_ _01949_ _01950_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__and2_1
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _08106_ _08107_ vssd1 vssd1 vccd1 vccd1 _08108_ sky130_fd_sc_hd__or2_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12675_ rbzero.debug_overlay.facingX\[-7\] rbzero.wall_tracer.rayAddendX\[1\] vssd1
+ vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__nor2_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17202_ _09782_ _09785_ vssd1 vssd1 vccd1 vccd1 _09786_ sky130_fd_sc_hd__xnor2_1
X_14414_ _07072_ _07148_ _07150_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__and3b_1
X_18182_ _01877_ _01882_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__xnor2_1
X_11626_ rbzero.tex_r1\[39\] rbzero.tex_r1\[38\] _04250_ vssd1 vssd1 vccd1 vccd1 _04405_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15394_ _07925_ _08037_ _08038_ vssd1 vssd1 vccd1 vccd1 _08039_ sky130_fd_sc_hd__a21o_2
X_17133_ _07706_ vssd1 vssd1 vccd1 vccd1 _09762_ sky130_fd_sc_hd__clkbuf_8
XFILLER_128_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14345_ _07015_ _07022_ _07081_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__a21oi_1
XFILLER_129_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11557_ _04128_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__buf_4
XFILLER_7_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10508_ rbzero.tex_r0\[35\] rbzero.tex_r0\[34\] _03580_ vssd1 vssd1 vccd1 vccd1 _03590_
+ sky130_fd_sc_hd__mux2_1
X_17064_ _05198_ _09703_ vssd1 vssd1 vccd1 vccd1 _09704_ sky130_fd_sc_hd__nand2_4
XFILLER_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11488_ _04258_ _04260_ _04267_ _04210_ _04242_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__a221o_1
XFILLER_144_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14276_ _07007_ _07012_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__xnor2_2
XFILLER_183_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16015_ _08111_ _08579_ vssd1 vssd1 vccd1 vccd1 _08660_ sky130_fd_sc_hd__nor2_1
X_10439_ rbzero.tex_r1\[1\] rbzero.tex_r1\[2\] _03549_ vssd1 vssd1 vccd1 vccd1 _03552_
+ sky130_fd_sc_hd__mux2_1
X_13227_ _05743_ _05874_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__o21a_1
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13158_ _05891_ _05892_ _05591_ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a2bb2o_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12109_ _04874_ _04876_ _04880_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__and3_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17966_ _01667_ _01668_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__nand2_1
X_13089_ _05795_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__clkbuf_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16917_ _09556_ _09557_ vssd1 vssd1 vccd1 vccd1 _09558_ sky130_fd_sc_hd__nand2_1
X_19705_ _03079_ vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17897_ _01593_ _01598_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__03305_ _03305_ vssd1 vssd1 vccd1 vccd1 clknet_0__03305_ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16848_ _08823_ _09028_ _09164_ _08329_ vssd1 vssd1 vccd1 vccd1 _09489_ sky130_fd_sc_hd__o22a_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19567_ _03034_ _03035_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__nor2_1
X_16779_ _09141_ _09420_ _08170_ vssd1 vssd1 vccd1 vccd1 _09421_ sky130_fd_sc_hd__a21oi_1
XFILLER_129_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18518_ _02102_ _02104_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__nor2_1
XFILLER_34_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19498_ rbzero.wall_tracer.rayAddendY\[6\] rbzero.wall_tracer.rayAddendY\[5\] _02905_
+ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__o21ai_1
XFILLER_55_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18449_ _02145_ _02146_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__nand2_1
XFILLER_22_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21460_ net381 _01229_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20411_ _02721_ _03322_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__and3_1
XFILLER_175_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21391_ net312 _01160_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20207__230 clknet_1_0__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__inv_2
XFILLER_72_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10790_ _03738_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ rbzero.wall_tracer.trackDistX\[9\] vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__inv_2
X_21658_ clknet_leaf_79_i_clk _01427_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11411_ gpout0.hpos\[2\] _04149_ _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__nand3b_1
XFILLER_123_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12391_ net41 _05139_ net34 net35 vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a211o_1
X_20609_ _03469_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xtop_ew_algofoogle_73 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_73/HI o_rgb[1] sky130_fd_sc_hd__conb_1
X_21589_ net130 _01358_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_84 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_84/HI o_rgb[16] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_95 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_95/HI zeros[5] sky130_fd_sc_hd__conb_1
XFILLER_181_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14130_ _06828_ _06864_ _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__a21o_1
X_11342_ _04092_ _04081_ _04089_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__nor3_1
XFILLER_193_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20253__272 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__inv_2
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11273_ _04048_ _04052_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__nand2_1
X_14061_ _06757_ _06797_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__xnor2_1
XFILLER_181_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13012_ _05695_ _05702_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__or3_1
XFILLER_121_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17820_ _10129_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__buf_2
XFILLER_121_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17751_ _10214_ _10230_ _10228_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a21o_1
XFILLER_181_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14963_ _07651_ vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__clkbuf_1
Xhold6 rbzero.wall_tracer.visualWallDist\[3\] vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16702_ _09210_ _09237_ _09343_ vssd1 vssd1 vccd1 vccd1 _09344_ sky130_fd_sc_hd__a21boi_1
XFILLER_43_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13914_ _06572_ _06627_ _06629_ _06650_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__o211a_1
X_17682_ _10245_ _10246_ vssd1 vssd1 vccd1 vccd1 _10247_ sky130_fd_sc_hd__xor2_2
XFILLER_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14894_ rbzero.wall_tracer.trackDistY\[-9\] rbzero.wall_tracer.trackDistX\[-9\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__mux2_1
XFILLER_130_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19421_ _02904_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__buf_2
XFILLER_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16633_ _08971_ vssd1 vssd1 vccd1 vccd1 _09276_ sky130_fd_sc_hd__clkbuf_4
XFILLER_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13845_ _06248_ _06581_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19352_ _02824_ _02837_ _02825_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__o21ai_1
X_16564_ _08549_ _08957_ _09204_ _09206_ vssd1 vssd1 vccd1 vccd1 _09207_ sky130_fd_sc_hd__a31o_4
X_13776_ _06406_ _06511_ _06512_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__a21bo_1
XFILLER_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10988_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _03762_ vssd1 vssd1 vccd1 vccd1 _03842_
+ sky130_fd_sc_hd__mux2_1
XFILLER_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18303_ _02001_ _02002_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__nor2_1
X_15515_ _08124_ vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__clkbuf_4
XFILLER_128_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12727_ _05473_ _05474_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__xnor2_2
X_19283_ _02796_ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__clkbuf_1
X_16495_ _08816_ _09138_ vssd1 vssd1 vccd1 vccd1 _09139_ sky130_fd_sc_hd__nor2_1
XFILLER_176_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18234_ _09661_ _09483_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__or2_2
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15446_ rbzero.wall_tracer.visualWallDist\[-1\] _08090_ _07951_ vssd1 vssd1 vccd1
+ vccd1 _08091_ sky130_fd_sc_hd__mux2_1
XFILLER_15_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12658_ rbzero.debug_overlay.playerY\[5\] _05407_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05408_ sky130_fd_sc_hd__mux2_1
XFILLER_50_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20336__347 clknet_1_1__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__inv_2
X_18165_ _09292_ _09695_ _09668_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a21o_1
X_11609_ rbzero.tex_r1\[55\] _04221_ _04222_ _04266_ vssd1 vssd1 vccd1 vccd1 _04388_
+ sky130_fd_sc_hd__a31o_1
XFILLER_191_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15377_ _08021_ vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__clkbuf_4
X_12589_ _05289_ _05295_ _05303_ _05301_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__a31o_1
XFILLER_102_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17116_ _05189_ vssd1 vssd1 vccd1 vccd1 _09753_ sky130_fd_sc_hd__buf_6
X_14328_ _07063_ _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18096_ _01796_ _01797_ _09817_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__o21a_1
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17047_ _09685_ _09686_ vssd1 vssd1 vccd1 vccd1 _09687_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14259_ _06724_ _06672_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__nor2_1
XFILLER_99_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19629__81 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__inv_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ rbzero.pov.spi_buffer\[31\] rbzero.pov.ready_buffer\[31\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02630_ sky130_fd_sc_hd__mux2_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17949_ _01650_ _01651_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__and2b_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20960_ clknet_leaf_7_i_clk _00729_ vssd1 vssd1 vccd1 vccd1 rbzero.otherx\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_66_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20081__117 clknet_1_0__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__inv_2
X_20891_ clknet_leaf_87_i_clk _00660_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21512_ net433 _01281_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21443_ net364 _01212_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21374_ net295 _01143_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11960_ rbzero.color_sky\[4\] rbzero.color_floor\[4\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04736_ sky130_fd_sc_hd__mux2_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10911_ rbzero.tex_b1\[35\] rbzero.tex_b1\[36\] _03795_ vssd1 vssd1 vccd1 vccd1 _03802_
+ sky130_fd_sc_hd__mux2_1
XFILLER_205_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ rbzero.tex_b0\[14\] _04291_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__and2_1
X_13630_ _06354_ _06366_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10842_ rbzero.tex_g0\[5\] rbzero.tex_g0\[4\] _03762_ vssd1 vssd1 vccd1 vccd1 _03766_
+ sky130_fd_sc_hd__mux2_1
XFILLER_198_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13561_ _06078_ _06161_ _06292_ _06297_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__o31a_1
X_10773_ rbzero.tex_g0\[38\] rbzero.tex_g0\[37\] _03729_ vssd1 vssd1 vccd1 vccd1 _03730_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15300_ _05207_ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__buf_6
XFILLER_40_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12512_ rbzero.wall_tracer.trackDistX\[-3\] vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__inv_2
XFILLER_197_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16280_ _08918_ vssd1 vssd1 vccd1 vccd1 _08925_ sky130_fd_sc_hd__inv_2
XFILLER_9_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13492_ _06175_ _06185_ _06228_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__a21oi_1
XFILLER_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15231_ _07821_ rbzero.wall_tracer.rayAddendX\[10\] vssd1 vssd1 vccd1 vccd1 _07881_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12443_ net71 rbzero.wall_tracer.state\[4\] _03480_ vssd1 vssd1 vccd1 vccd1 _05200_
+ sky130_fd_sc_hd__and3_1
XFILLER_154_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15162_ _07785_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _07817_
+ sky130_fd_sc_hd__or2_1
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12374_ net33 vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__inv_2
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14113_ _06691_ _06849_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__xnor2_1
XFILLER_153_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11325_ _04103_ _04104_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15093_ _07738_ _07752_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__or2_1
X_19970_ rbzero.pov.ready_buffer\[43\] _03240_ _03243_ rbzero.debug_overlay.facingX\[10\]
+ _03244_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__o221a_1
XFILLER_158_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11256_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__buf_4
X_18921_ rbzero.spi_registers.spi_counter\[4\] _02583_ vssd1 vssd1 vccd1 vccd1 _02587_
+ sky130_fd_sc_hd__or2_1
X_14044_ _06774_ _06775_ _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__and3_1
XFILLER_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18852_ _02524_ _02525_ _02526_ _05531_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a31o_1
X_11187_ _03974_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__nand2_1
XFILLER_95_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17803_ _01505_ _01506_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__xor2_2
XFILLER_132_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18783_ _02465_ _02466_ _02467_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__o21a_1
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15995_ _08633_ _08632_ vssd1 vssd1 vccd1 vccd1 _08640_ sky130_fd_sc_hd__xor2_1
XFILLER_48_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17734_ _09812_ _10181_ _10182_ _05414_ _01438_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__o311a_1
X_14946_ rbzero.wall_tracer.trackDistY\[7\] rbzero.wall_tracer.trackDistX\[7\] _05278_
+ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__mux2_1
XFILLER_76_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17665_ _10228_ _10229_ vssd1 vssd1 vccd1 vccd1 _10230_ sky130_fd_sc_hd__nor2_1
X_14877_ _07590_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16616_ _09256_ _09258_ vssd1 vssd1 vccd1 vccd1 _09259_ sky130_fd_sc_hd__nor2_1
X_19404_ _02883_ _02888_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__nand2_1
X_13828_ _06268_ _06235_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__or2b_1
XFILLER_91_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17596_ _09918_ _10018_ _10161_ vssd1 vssd1 vccd1 vccd1 _10162_ sky130_fd_sc_hd__a21boi_1
XFILLER_165_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16547_ _09053_ _09189_ _09190_ vssd1 vssd1 vccd1 vccd1 _09191_ sky130_fd_sc_hd__a21oi_2
X_19335_ _02824_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__and2b_1
X_13759_ _06461_ _06458_ _06465_ _06495_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__a211o_1
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19266_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_floor\[3\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__mux2_1
X_16478_ _08383_ _07959_ vssd1 vssd1 vccd1 vccd1 _09122_ sky130_fd_sc_hd__nor2_1
X_18217_ _01688_ _01690_ _01816_ _01814_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__a31o_1
XFILLER_176_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15429_ _05206_ _08068_ _08072_ _08073_ vssd1 vssd1 vccd1 vccd1 _08074_ sky130_fd_sc_hd__a22o_2
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19197_ rbzero.spi_registers.new_sky\[2\] rbzero.spi_registers.got_new_sky _02711_
+ _02741_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a31o_1
XFILLER_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18148_ _01716_ _01725_ _01724_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__o21ba_1
XFILLER_157_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18079_ _01697_ _01780_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21090_ net180 _00859_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20041_ _04886_ _04990_ _03275_ _03911_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__a31o_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20943_ clknet_leaf_10_i_clk _00712_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ clknet_leaf_95_i_clk _00643_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20319__331 clknet_1_0__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__inv_2
XFILLER_33_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21426_ net347 _01195_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21357_ net278 _01126_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11110_ rbzero.tex_b0\[5\] rbzero.tex_b0\[4\] _03898_ vssd1 vssd1 vccd1 vccd1 _03906_
+ sky130_fd_sc_hd__mux2_1
XFILLER_107_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12090_ _04851_ _04856_ _04861_ _04850_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a22o_1
X_21288_ clknet_leaf_37_i_clk _01057_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11041_ rbzero.tex_b0\[38\] rbzero.tex_b0\[37\] _03865_ vssd1 vssd1 vccd1 vccd1 _03870_
+ sky130_fd_sc_hd__mux2_1
X_19608__62 clknet_1_1__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__inv_2
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ rbzero.wall_tracer.stepDistY\[-6\] _07461_ vssd1 vssd1 vccd1 vccd1 _07531_
+ sky130_fd_sc_hd__nor2_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20365__373 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__inv_2
X_19623__76 clknet_1_1__leaf__03042_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__inv_2
XFILLER_64_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15780_ _08424_ vssd1 vssd1 vccd1 vccd1 _08425_ sky130_fd_sc_hd__clkbuf_2
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12992_ _05728_ _05645_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__nand2_1
XFILLER_188_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20064__101 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__inv_2
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14731_ _07466_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__clkbuf_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11943_ _04717_ _04718_ _04329_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__mux2_1
XFILLER_206_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17450_ _09657_ _09725_ _10016_ vssd1 vssd1 vccd1 vccd1 _10017_ sky130_fd_sc_hd__a21o_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _05892_ _07395_ _07398_ _07375_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__o211a_1
X_11874_ _04649_ _04650_ _04224_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__mux2_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16401_ _08367_ _09026_ _09044_ vssd1 vssd1 vccd1 vccd1 _09046_ sky130_fd_sc_hd__nand3_2
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13613_ _06345_ _06346_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__xnor2_1
X_17381_ _09521_ _09525_ _09645_ vssd1 vssd1 vccd1 vccd1 _09948_ sky130_fd_sc_hd__a21oi_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10825_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _03751_ vssd1 vssd1 vccd1 vccd1 _03757_
+ sky130_fd_sc_hd__mux2_1
X_14593_ _07213_ _07328_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__nand2_1
XFILLER_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19120_ _02694_ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__clkbuf_1
X_16332_ _07602_ _08230_ _08147_ _08225_ vssd1 vssd1 vccd1 vccd1 _08977_ sky130_fd_sc_hd__or4b_2
XFILLER_185_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13544_ _06132_ _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__xor2_2
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10756_ rbzero.tex_g0\[46\] rbzero.tex_g0\[45\] _03718_ vssd1 vssd1 vccd1 vccd1 _03721_
+ sky130_fd_sc_hd__mux2_1
XFILLER_201_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19051_ _02657_ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__clkbuf_1
X_16263_ _08897_ _08907_ vssd1 vssd1 vccd1 vccd1 _08908_ sky130_fd_sc_hd__xor2_1
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13475_ _05910_ _06176_ _06085_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__and3_1
X_10687_ _03684_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__clkbuf_1
X_18002_ _09249_ _09703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__and2_1
X_15214_ _07843_ _07845_ _07864_ _07676_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__a31o_1
XFILLER_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12426_ _03480_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__buf_4
XFILLER_199_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16194_ _08793_ _08838_ vssd1 vssd1 vccd1 vccd1 _08839_ sky130_fd_sc_hd__or2_1
XFILLER_127_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15145_ _07742_ rbzero.debug_overlay.vplaneX\[-4\] vssd1 vssd1 vccd1 vccd1 _07801_
+ sky130_fd_sc_hd__and2_1
X_12357_ net49 _05084_ _05107_ net50 vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__a22o_1
XFILLER_153_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ _04084_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__or2_1
X_15076_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__nand2_1
X_19953_ rbzero.pov.ready_buffer\[34\] _03240_ _03243_ rbzero.debug_overlay.facingX\[-8\]
+ _03209_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__o221a_1
X_12288_ net39 _05046_ _05049_ net40 vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a22o_1
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18904_ _02557_ _02573_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__and2_1
X_14027_ _06704_ _06761_ _06763_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__or3_1
X_11239_ gpout0.hpos\[2\] gpout0.hpos\[1\] gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1
+ _04023_ sky130_fd_sc_hd__and3_2
X_19884_ _03189_ _03191_ _02714_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__o21a_1
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18835_ _02510_ _02511_ _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a21oi_1
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15978_ _07912_ _08328_ _08040_ vssd1 vssd1 vccd1 vccd1 _08623_ sky130_fd_sc_hd__or3b_2
X_18766_ _02443_ _02445_ _02444_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a21boi_1
XFILLER_48_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17717_ _10152_ _10154_ vssd1 vssd1 vccd1 vccd1 _10282_ sky130_fd_sc_hd__nor2_1
X_14929_ rbzero.wall_tracer.visualWallDist\[1\] _07618_ vssd1 vssd1 vccd1 vccd1 _07629_
+ sky130_fd_sc_hd__or2_1
X_18697_ _02391_ _02392_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__xnor2_1
XFILLER_63_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17648_ _10211_ _10212_ vssd1 vssd1 vccd1 vccd1 _10213_ sky130_fd_sc_hd__nor2_1
XFILLER_1_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17579_ _10127_ _10136_ _10142_ _10144_ vssd1 vssd1 vccd1 vccd1 _10145_ sky130_fd_sc_hd__o22a_1
XFILLER_177_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19318_ _02815_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20590_ rbzero.debug_overlay.vplaneY\[-9\] rbzero.wall_tracer.rayAddendY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__or2_1
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20193__218 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__inv_2
XFILLER_164_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19249_ _02777_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21211_ clknet_leaf_26_i_clk _00980_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21142_ clknet_leaf_97_i_clk _00911_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21073_ net163 _00842_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20024_ _04992_ _03267_ _03268_ _03209_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__o211a_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ clknet_leaf_26_i_clk _00695_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20857_ clknet_leaf_1_i_clk _00626_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10610_ _03643_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__clkbuf_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11590_ rbzero.tex_r1\[30\] _04350_ _04265_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__a21o_1
X_20788_ clknet_leaf_47_i_clk _00557_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _03607_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ _05993_ _05996_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__or2b_1
X_10472_ _03571_ vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12211_ _04960_ _04961_ _04963_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__and3_1
XFILLER_109_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21409_ net330 _01178_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[52\] sky130_fd_sc_hd__dfxtp_1
X_13191_ _05743_ _05754_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__nor2_2
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _04910_ _04738_ net12 net11 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__o211a_1
XFILLER_155_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12073_ _04840_ net66 _04844_ net6 vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__a211o_1
X_16950_ _09345_ _09590_ vssd1 vssd1 vccd1 vccd1 _09591_ sky130_fd_sc_hd__xor2_1
XFILLER_81_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15901_ _08509_ _08544_ _08545_ vssd1 vssd1 vccd1 vccd1 _08546_ sky130_fd_sc_hd__a21oi_2
X_11024_ rbzero.tex_b0\[46\] rbzero.tex_b0\[45\] _03854_ vssd1 vssd1 vccd1 vccd1 _03861_
+ sky130_fd_sc_hd__mux2_1
X_16881_ _07994_ vssd1 vssd1 vccd1 vccd1 _09522_ sky130_fd_sc_hd__buf_2
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15832_ _08473_ _08474_ _08476_ vssd1 vssd1 vccd1 vccd1 _08477_ sky130_fd_sc_hd__a21bo_1
X_18620_ rbzero.wall_tracer.trackDistX\[10\] rbzero.wall_tracer.stepDistX\[10\] vssd1
+ vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__or2_1
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _02236_ _02247_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__xnor2_1
X_15763_ _08406_ _08407_ vssd1 vssd1 vccd1 vccd1 _08408_ sky130_fd_sc_hd__nand2_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12975_ _05594_ _05596_ _05598_ _05584_ _05628_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__o41a_2
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17502_ _10057_ _10066_ vssd1 vssd1 vccd1 vccd1 _10068_ sky130_fd_sc_hd__or2_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14714_ _07348_ _07353_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__nand2_1
X_18482_ _02176_ _02178_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__nand2_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ rbzero.tex_b0\[61\] rbzero.tex_b0\[60\] _04263_ vssd1 vssd1 vccd1 vccd1 _04702_
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15694_ _08084_ _07964_ _07965_ vssd1 vssd1 vccd1 vccd1 _08339_ sky130_fd_sc_hd__or3_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _09700_ _09997_ _09998_ _09999_ vssd1 vssd1 vccd1 vccd1 _10000_ sky130_fd_sc_hd__o2bb2a_2
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14645_ _05931_ _07381_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__nor2_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ rbzero.tex_g1\[11\] _04327_ _04328_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__and3_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17364_ _09929_ _09930_ vssd1 vssd1 vccd1 vccd1 _09931_ sky130_fd_sc_hd__xor2_1
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10808_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _03740_ vssd1 vssd1 vccd1 vccd1 _03748_
+ sky130_fd_sc_hd__mux2_1
X_14576_ _07095_ _07035_ _07043_ _07098_ _07312_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__a221o_1
XFILLER_207_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11788_ rbzero.tex_g0\[51\] rbzero.tex_g0\[50\] _04262_ vssd1 vssd1 vccd1 vccd1 _04566_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16315_ _08008_ _08204_ vssd1 vssd1 vccd1 vccd1 _08960_ sky130_fd_sc_hd__or2_1
X_19103_ rbzero.spi_registers.spi_buffer\[7\] rbzero.spi_registers.spi_buffer\[6\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__mux2_1
XFILLER_203_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13527_ _06256_ _06257_ _06262_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__or3_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10739_ _03711_ vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__clkbuf_1
X_17295_ _09864_ _09865_ _09866_ vssd1 vssd1 vccd1 vccd1 _09867_ sky130_fd_sc_hd__and3_1
XFILLER_185_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19034_ _02648_ vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__clkbuf_1
X_16246_ _08879_ _08883_ _08890_ vssd1 vssd1 vccd1 vccd1 _08891_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _06191_ _06189_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__or2b_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12409_ _05171_ _05175_ net36 vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__or3b_1
X_16177_ _08112_ _08328_ _08747_ vssd1 vssd1 vccd1 vccd1 _08822_ sky130_fd_sc_hd__or3_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13389_ _06121_ _06124_ _06125_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__and3_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15128_ rbzero.debug_overlay.vplaneX\[10\] vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15059_ rbzero.debug_overlay.vplaneX\[-2\] rbzero.wall_tracer.rayAddendX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__or2_1
X_19936_ _02820_ _03227_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__nor2_1
XFILLER_130_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19867_ _03176_ _03177_ _02822_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18818_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.stepDistY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__or2_1
XFILLER_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19798_ rbzero.pov.spi_buffer\[72\] rbzero.pov.spi_buffer\[73\] _03047_ vssd1 vssd1
+ vccd1 vccd1 _03128_ sky130_fd_sc_hd__mux2_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18749_ _02435_ _02436_ _02437_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__nor3_1
XFILLER_97_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19602__57 clknet_1_1__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__03298_ clknet_0__03298_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03298_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20711_ clknet_leaf_72_i_clk _00002_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20201__225 clknet_1_1__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__inv_2
X_20642_ clknet_leaf_64_i_clk _00426_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20573_ _03447_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_165_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_opt_1_0_i_clk clknet_3_0_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_1_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_149_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21125_ clknet_leaf_95_i_clk _00894_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_121_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21056_ clknet_leaf_0_i_clk _00825_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20007_ _03020_ _03019_ _03025_ rbzero.pov.spi_done vssd1 vssd1 vccd1 vccd1 _03255_
+ sky130_fd_sc_hd__a31o_1
XFILLER_47_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _03924_ _05503_ _05499_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__o21ai_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _04481_ _04489_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__nand2_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ clknet_leaf_92_i_clk _00678_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _05421_ _05430_ _05433_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__a31o_1
XFILLER_187_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _07137_ _07045_ _07165_ _07166_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_202_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11642_ _04414_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__inv_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20176__202 clknet_1_1__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__inv_2
XFILLER_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14361_ _07095_ _07097_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__xnor2_1
X_11573_ rbzero.tex_r1\[1\] rbzero.tex_r1\[0\] _04342_ vssd1 vssd1 vccd1 vccd1 _04352_
+ sky130_fd_sc_hd__mux2_1
XFILLER_126_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16100_ _08519_ _08075_ _08674_ _08377_ vssd1 vssd1 vccd1 vccd1 _08745_ sky130_fd_sc_hd__o22ai_2
Xinput18 i_gpout2_sel[4] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_8
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13312_ _06022_ _06038_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__nand2_1
X_10524_ _03598_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__clkbuf_1
X_17080_ _09550_ _09574_ _09719_ vssd1 vssd1 vccd1 vccd1 _09720_ sky130_fd_sc_hd__a21oi_2
Xinput29 i_gpout4_sel[3] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_6
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14292_ _06737_ _06817_ _07028_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__a21boi_2
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16031_ _07980_ _07964_ _07965_ vssd1 vssd1 vccd1 vccd1 _08676_ sky130_fd_sc_hd__or3_1
X_13243_ _05979_ _05899_ _05846_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__o21ai_2
XFILLER_109_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10455_ _03562_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13174_ _05867_ _05783_ _05792_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__mux2_1
XFILLER_163_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10386_ rbzero.tex_r1\[26\] rbzero.tex_r1\[27\] _03516_ vssd1 vssd1 vccd1 vccd1 _03524_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12125_ _04852_ clknet_1_1__leaf__04835_ _04855_ gpout0.clk_div\[1\] _04838_ vssd1
+ vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__a221o_2
XFILLER_2_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17982_ _01660_ _01662_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__or2_1
X_19721_ rbzero.pov.spi_buffer\[35\] rbzero.pov.spi_buffer\[36\] _03081_ vssd1 vssd1
+ vccd1 vccd1 _03088_ sky130_fd_sc_hd__mux2_1
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12056_ _04819_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__nor2_1
X_16933_ _09571_ _09573_ vssd1 vssd1 vccd1 vccd1 _09574_ sky130_fd_sc_hd__xnor2_2
XFILLER_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03321_ _03321_ vssd1 vssd1 vccd1 vccd1 clknet_0__03321_ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ rbzero.tex_b0\[54\] rbzero.tex_b0\[53\] _03843_ vssd1 vssd1 vccd1 vccd1 _03852_
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19652_ rbzero.pov.spi_buffer\[2\] rbzero.pov.spi_buffer\[3\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03052_ sky130_fd_sc_hd__mux2_1
XFILLER_38_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16864_ _09501_ _09504_ vssd1 vssd1 vccd1 vccd1 _09505_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18603_ _02208_ _02299_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__xnor2_1
XFILLER_168_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15815_ _08441_ _08459_ vssd1 vssd1 vccd1 vccd1 _08460_ sky130_fd_sc_hd__xor2_1
XFILLER_19_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16795_ _09290_ _09291_ vssd1 vssd1 vccd1 vccd1 _09437_ sky130_fd_sc_hd__nand2_1
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18534_ _02229_ _02230_ _02231_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a21oi_1
X_15746_ _08373_ _08390_ vssd1 vssd1 vccd1 vccd1 _08391_ sky130_fd_sc_hd__xnor2_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ _05674_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__buf_2
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11909_ rbzero.tex_b0\[17\] rbzero.tex_b0\[16\] _04271_ vssd1 vssd1 vccd1 vccd1 _04685_
+ sky130_fd_sc_hd__mux2_1
X_18465_ _02161_ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__xor2_1
X_15677_ _08321_ _08286_ vssd1 vssd1 vccd1 vccd1 _08322_ sky130_fd_sc_hd__xnor2_1
XFILLER_34_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12889_ _04001_ _05456_ _05624_ _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a22oi_4
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17416_ _09114_ _09417_ vssd1 vssd1 vccd1 vccd1 _09983_ sky130_fd_sc_hd__nor2_1
X_14628_ _07363_ _07364_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__xnor2_1
XFILLER_178_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18396_ _01952_ _01959_ _02094_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17347_ _09912_ _09913_ vssd1 vssd1 vccd1 vccd1 _09914_ sky130_fd_sc_hd__or2_1
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14559_ _07289_ _07290_ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__or2_1
XFILLER_140_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _09812_ _09849_ _09850_ _09851_ vssd1 vssd1 vccd1 vccd1 _09852_ sky130_fd_sc_hd__o31ai_1
XFILLER_173_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16229_ _08872_ _08491_ _08579_ _08873_ vssd1 vssd1 vccd1 vccd1 _08874_ sky130_fd_sc_hd__o22a_1
X_19017_ rbzero.pov.spi_buffer\[40\] rbzero.pov.ready_buffer\[40\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02640_ sky130_fd_sc_hd__mux2_1
XFILLER_174_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19919_ rbzero.debug_overlay.playerY\[0\] _08030_ vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__nand2_1
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03310_ clknet_0__03310_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03310_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_178_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20625_ clknet_leaf_16_i_clk _00409_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f2 sky130_fd_sc_hd__dfxtp_2
XFILLER_193_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20556_ _07695_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__buf_4
XFILLER_192_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20487_ _03383_ _03384_ _03385_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__and3_1
XFILLER_118_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20171__198 clknet_1_1__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__inv_2
XFILLER_161_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21108_ net198 _00877_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13930_ _06603_ _06612_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__xnor2_4
XFILLER_75_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21039_ clknet_leaf_74_i_clk _00808_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_93_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13861_ _06277_ _06563_ _06597_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__o21bai_4
X_15600_ _08243_ _08244_ vssd1 vssd1 vccd1 vccd1 _08245_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12812_ rbzero.wall_tracer.mapY\[9\] _05404_ _05550_ vssd1 vssd1 vccd1 vccd1 _05552_
+ sky130_fd_sc_hd__o21a_1
X_16580_ _09170_ _09172_ _09169_ vssd1 vssd1 vccd1 vccd1 _09223_ sky130_fd_sc_hd__a21bo_1
XFILLER_90_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13792_ _06527_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__xnor2_1
XFILLER_16_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15531_ _08148_ rbzero.wall_tracer.stepDistY\[1\] _07990_ vssd1 vssd1 vccd1 vccd1
+ _08176_ sky130_fd_sc_hd__o21a_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _05459_ _05484_ _05488_ _05490_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__and4b_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18250_ _01938_ _01948_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_91_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _08086_ _08087_ _08105_ vssd1 vssd1 vccd1 vccd1 _08107_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ rbzero.debug_overlay.facingX\[-6\] rbzero.wall_tracer.rayAddendX\[2\] vssd1
+ vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__nor2_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _09783_ _09784_ vssd1 vssd1 vccd1 vccd1 _09785_ sky130_fd_sc_hd__or2_1
X_14413_ _06760_ _07117_ _07149_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__or3b_1
X_18181_ _01756_ _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__xnor2_1
XFILLER_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ _04266_ _04403_ _04229_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__o21a_1
X_15393_ _07904_ rbzero.wall_tracer.stepDistY\[-9\] _05206_ vssd1 vssd1 vccd1 vccd1
+ _08038_ sky130_fd_sc_hd__a21o_1
XFILLER_128_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17132_ _09760_ _09761_ _09748_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14344_ _07020_ _07021_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__and2_1
XFILLER_155_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11556_ rbzero.tex_r1\[11\] _04327_ _04328_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__and3_1
XFILLER_183_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10507_ _03589_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__clkbuf_1
X_17063_ _03953_ _09283_ vssd1 vssd1 vccd1 vccd1 _09703_ sky130_fd_sc_hd__nor2_4
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14275_ _07008_ _07011_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__xnor2_1
X_11487_ _04261_ _04264_ _04266_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__mux2_1
X_16014_ _08573_ _08575_ vssd1 vssd1 vccd1 vccd1 _08659_ sky130_fd_sc_hd__xnor2_1
XFILLER_100_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13226_ _05928_ _05901_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__nor2_1
XFILLER_171_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ _03551_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _05743_ _05826_ _05893_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__and3_1
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10369_ rbzero.tex_r1\[34\] rbzero.tex_r1\[35\] _03505_ vssd1 vssd1 vccd1 vccd1 _03515_
+ sky130_fd_sc_hd__mux2_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20230__251 clknet_1_0__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__inv_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12108_ _04877_ _04878_ _04879_ _04869_ net7 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__o221a_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17965_ _01664_ _01666_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__nand2_1
X_13088_ _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__buf_4
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19704_ rbzero.pov.spi_buffer\[27\] rbzero.pov.spi_buffer\[28\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03079_ sky130_fd_sc_hd__mux2_1
X_12039_ _04022_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__buf_2
X_16916_ _08873_ _09540_ _09555_ _08872_ vssd1 vssd1 vccd1 vccd1 _09557_ sky130_fd_sc_hd__o22ai_1
XFILLER_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17896_ _01593_ _01598_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__and2_1
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03304_ _03304_ vssd1 vssd1 vccd1 vccd1 clknet_0__03304_ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_16847_ _08054_ _09216_ vssd1 vssd1 vccd1 vccd1 _09488_ sky130_fd_sc_hd__nor2_1
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20148__178 clknet_1_1__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__inv_2
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19566_ rbzero.pov.spi_counter\[5\] _03031_ _03020_ vssd1 vssd1 vccd1 vccd1 _03035_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_53_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16778_ _05210_ rbzero.wall_tracer.stepDistX\[6\] vssd1 vssd1 vccd1 vccd1 _09420_
+ sky130_fd_sc_hd__nand2_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18517_ _02204_ _02214_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__xnor2_2
X_15729_ _08188_ _08238_ vssd1 vssd1 vccd1 vccd1 _08374_ sky130_fd_sc_hd__nor2_1
X_19497_ _02950_ _02951_ _02968_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_59_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18448_ _10238_ _09292_ _09991_ _01737_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__o22ai_1
XFILLER_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18379_ _02075_ _02077_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__or2_1
XFILLER_144_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20410_ gpout5.clk_div\[1\] gpout5.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__or2_1
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21390_ net311 _01159_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20313__326 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__inv_2
XFILLER_162_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20272_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__buf_1
XFILLER_161_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21657_ clknet_leaf_91_i_clk _01426_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11410_ _04147_ _04148_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__or2_1
XFILLER_123_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20608_ _02721_ _03467_ _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__and3_1
XFILLER_137_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ net39 _05144_ _05156_ _05153_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a211o_1
XFILLER_193_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21588_ net509 _01357_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xtop_ew_algofoogle_74 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_74/HI o_rgb[2] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_85 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_85/HI o_rgb[17] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_96 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_96/HI zeros[6] sky130_fd_sc_hd__conb_1
XFILLER_123_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11341_ _04100_ _04114_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__or3_4
XFILLER_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20539_ rbzero.traced_texa\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _03430_
+ sky130_fd_sc_hd__or2_1
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14060_ _06784_ _06796_ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__xnor2_1
XFILLER_152_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11272_ rbzero.traced_texVinit\[9\] rbzero.texV\[9\] vssd1 vssd1 vccd1 vccd1 _04052_
+ sky130_fd_sc_hd__or2_1
XFILLER_118_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20288__303 clknet_1_0__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__inv_2
X_13011_ _05691_ _05744_ _05682_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__or3_1
XFILLER_165_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17750_ _10189_ _01453_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14962_ rbzero.wall_tracer.stepDistX\[-12\] _07460_ _07650_ vssd1 vssd1 vccd1 vccd1
+ _07651_ sky130_fd_sc_hd__mux2_1
XFILLER_43_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16701_ _09238_ _09209_ vssd1 vssd1 vccd1 vccd1 _09343_ sky130_fd_sc_hd__or2b_1
XFILLER_48_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13913_ _06632_ _06649_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__xnor2_1
X_17681_ _09276_ _09674_ vssd1 vssd1 vccd1 vccd1 _10246_ sky130_fd_sc_hd__nor2_1
XFILLER_43_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14893_ _07591_ _07600_ _07603_ _04039_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__o211a_1
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19420_ rbzero.debug_overlay.vplaneY\[10\] vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__clkbuf_4
X_16632_ _09268_ _09274_ vssd1 vssd1 vccd1 vccd1 _09275_ sky130_fd_sc_hd__xnor2_1
XFILLER_130_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13844_ _06579_ _06580_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__and2_1
XFILLER_207_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19351_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__and2_1
X_16563_ _09089_ _09205_ _09192_ vssd1 vssd1 vccd1 vccd1 _09206_ sky130_fd_sc_hd__a21boi_1
XFILLER_16_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13775_ _06061_ _06009_ _06510_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__o21bai_1
X_10987_ _03841_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18302_ _01890_ _01892_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__and2_1
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15514_ _08158_ vssd1 vssd1 vccd1 vccd1 _08159_ sky130_fd_sc_hd__clkbuf_4
X_12726_ _05423_ _05426_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__and2b_1
X_16494_ _08230_ rbzero.wall_tracer.stepDistY\[7\] _08235_ _09137_ vssd1 vssd1 vccd1
+ vccd1 _09138_ sky130_fd_sc_hd__a22oi_4
X_19282_ rbzero.spi_registers.spi_buffer\[3\] rbzero.spi_registers.new_leak\[3\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__mux2_1
XFILLER_188_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18233_ _09661_ _09480_ _09484_ _01462_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__o22ai_1
XFILLER_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15445_ _08089_ rbzero.debug_overlay.playerY\[-1\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _08090_ sky130_fd_sc_hd__mux2_2
X_12657_ _05405_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ rbzero.tex_r1\[54\] _04273_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__and2_1
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18164_ _01863_ _01864_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__and2_1
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15376_ _08019_ _08020_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__or2_1
XFILLER_156_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12588_ _05332_ _05341_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__and2_1
X_17115_ _09752_ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__clkbuf_1
X_14327_ _06680_ _06739_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__or2_1
XFILLER_184_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11539_ gpout0.hpos\[0\] _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__nand2_1
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18095_ _01793_ _01794_ _01795_ _09863_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__a31o_1
XFILLER_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17046_ _08237_ _09279_ _08283_ vssd1 vssd1 vccd1 vccd1 _09686_ sky130_fd_sc_hd__a21oi_2
X_14258_ _06882_ _06883_ _06994_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__nor3_4
XFILLER_99_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ _05852_ _05853_ _05855_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__a21oi_2
X_14189_ _05984_ _06671_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__nor2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _02629_ vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__clkbuf_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17948_ _01647_ _01648_ _01649_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a21o_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20403__28 clknet_1_0__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__inv_2
X_17879_ _07974_ _09164_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__or2_1
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20890_ clknet_leaf_86_i_clk _00659_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19549_ rbzero.pov.spi_counter\[1\] rbzero.pov.spi_counter\[0\] _03019_ vssd1 vssd1
+ vccd1 vccd1 _03022_ sky130_fd_sc_hd__and3_1
XFILLER_81_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19572__29 clknet_1_1__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__inv_2
XFILLER_55_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21511_ net432 _01280_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21442_ net363 _01211_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21373_ net294 _01142_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10910_ _03801_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__clkbuf_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _04666_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkinv_4
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10841_ _03765_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13560_ _06293_ _06296_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__nand2_1
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10772_ _03717_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__clkbuf_4
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12511_ _05263_ rbzero.wall_tracer.trackDistY\[-4\] _05265_ vssd1 vssd1 vccd1 vccd1
+ _05266_ sky130_fd_sc_hd__a21o_1
XFILLER_160_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13491_ _06173_ _06186_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__nor2_1
X_15230_ _07879_ vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__inv_2
XFILLER_185_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _05199_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15161_ _07785_ rbzero.wall_tracer.rayAddendX\[5\] vssd1 vssd1 vccd1 vccd1 _07816_
+ sky130_fd_sc_hd__nand2_1
X_12373_ net34 net64 _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__nor3b_1
XFILLER_138_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14112_ _06681_ _06688_ _06693_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__a21oi_1
XFILLER_10_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ rbzero.texV\[7\] _04058_ _04057_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__a21boi_1
XFILLER_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15092_ _07750_ _07751_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__and2_1
XFILLER_10_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18920_ rbzero.spi_registers.spi_counter\[4\] _02583_ vssd1 vssd1 vccd1 vccd1 _02586_
+ sky130_fd_sc_hd__nand2_1
X_14043_ _06777_ _06778_ _06779_ _06773_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__a22o_1
X_11255_ _04020_ _04026_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__and2_1
XFILLER_107_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18851_ _02524_ _02525_ _02526_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a21oi_1
X_11186_ rbzero.map_rom.f2 _03933_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__or2_1
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17802_ _09674_ _09417_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__nor2_1
XFILLER_132_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18782_ _02457_ _02459_ _02458_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__a21boi_1
X_15994_ _08589_ _08598_ vssd1 vssd1 vccd1 vccd1 _08639_ sky130_fd_sc_hd__xnor2_1
XFILLER_134_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17733_ _09812_ _10297_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__nand2_1
X_14945_ _07621_ _07638_ _07639_ _07620_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__o211a_1
XFILLER_78_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17664_ _10225_ _10227_ vssd1 vssd1 vccd1 vccd1 _10229_ sky130_fd_sc_hd__and2_1
X_14876_ rbzero.wall_tracer.stepDistY\[11\] _07589_ _05188_ vssd1 vssd1 vccd1 vccd1
+ _07590_ sky130_fd_sc_hd__mux2_1
X_20342__352 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__inv_2
XFILLER_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19403_ _02883_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__or2_1
XFILLER_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16615_ _07932_ _09103_ _09100_ _09257_ vssd1 vssd1 vccd1 vccd1 _09258_ sky130_fd_sc_hd__o31a_1
XFILLER_90_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13827_ _06232_ _06275_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__and2_1
X_17595_ _10015_ _10017_ vssd1 vssd1 vccd1 vccd1 _10161_ sky130_fd_sc_hd__or2b_1
XFILLER_91_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19334_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__nand2_1
X_16546_ _09050_ _09052_ vssd1 vssd1 vccd1 vccd1 _09190_ sky130_fd_sc_hd__nor2_1
X_13758_ _06490_ _06493_ _06494_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12709_ _05444_ _05443_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__or2b_1
X_19265_ _02786_ vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__clkbuf_1
X_16477_ _08963_ _09119_ _09120_ vssd1 vssd1 vccd1 vccd1 _09121_ sky130_fd_sc_hd__a21bo_1
X_13689_ _06379_ _06421_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__xnor2_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18216_ _01900_ _01804_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__or2b_1
X_15428_ rbzero.wall_tracer.visualWallDist\[-3\] _04013_ _05206_ vssd1 vssd1 vccd1
+ vccd1 _08073_ sky130_fd_sc_hd__a21oi_1
XFILLER_176_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19196_ _02744_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_89_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18147_ _01839_ _01847_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__xnor2_1
XFILLER_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15359_ _07905_ _08003_ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__and2_1
XFILLER_144_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18078_ _01777_ _01779_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__xor2_1
XFILLER_7_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17029_ _08178_ _09668_ vssd1 vssd1 vccd1 vccd1 _09669_ sky130_fd_sc_hd__nor2_2
XFILLER_172_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20040_ _04990_ _03275_ _03279_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__o21a_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_864 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ clknet_leaf_2_i_clk _00711_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_113_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ clknet_leaf_95_i_clk _00642_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21425_ net346 _01194_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21356_ net277 _01125_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21287_ clknet_leaf_35_i_clk _01056_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[5\] sky130_fd_sc_hd__dfxtp_4
XFILLER_150_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11040_ _03869_ vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__clkbuf_1
X_20238_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__buf_1
XFILLER_76_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _05609_ _05641_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__xnor2_1
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14730_ rbzero.wall_tracer.stepDistY\[-11\] _07465_ _07461_ vssd1 vssd1 vccd1 vccd1
+ _07466_ sky130_fd_sc_hd__mux2_1
X_11942_ rbzero.tex_b0\[41\] rbzero.tex_b0\[40\] _04342_ vssd1 vssd1 vccd1 vccd1 _04718_
+ sky130_fd_sc_hd__mux2_1
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20394__19 clknet_1_1__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__inv_2
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _05741_ _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__or2_1
X_11873_ rbzero.tex_g1\[23\] rbzero.tex_g1\[22\] _04211_ vssd1 vssd1 vccd1 vccd1 _04650_
+ sky130_fd_sc_hd__mux2_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16400_ _08367_ _09026_ _09044_ vssd1 vssd1 vccd1 vccd1 _09045_ sky130_fd_sc_hd__a21o_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13612_ _06348_ _06326_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__xnor2_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10824_ _03756_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__clkbuf_1
X_17380_ _09939_ _09946_ vssd1 vssd1 vccd1 vccd1 _09947_ sky130_fd_sc_hd__xnor2_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _07213_ _07328_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__nor2_1
XFILLER_77_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16331_ _08974_ _08975_ vssd1 vssd1 vccd1 vccd1 _08976_ sky130_fd_sc_hd__xnor2_2
XFILLER_125_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13543_ _06135_ _06133_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nor2_1
X_10755_ _03720_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16262_ _08905_ _08906_ vssd1 vssd1 vccd1 vccd1 _08907_ sky130_fd_sc_hd__and2b_1
X_19050_ rbzero.pov.spi_buffer\[56\] rbzero.pov.ready_buffer\[56\] _02649_ vssd1 vssd1
+ vccd1 vccd1 _02657_ sky130_fd_sc_hd__mux2_1
XFILLER_200_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13474_ _06157_ _06166_ _06210_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__a21bo_1
XFILLER_199_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10686_ rbzero.tex_g1\[14\] rbzero.tex_g1\[15\] _03680_ vssd1 vssd1 vccd1 vccd1 _03684_
+ sky130_fd_sc_hd__mux2_1
X_18001_ _01701_ _01702_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__or2_1
XFILLER_185_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15213_ _07843_ _07845_ _07864_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__a21oi_1
X_12425_ _04032_ _03914_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__nor2_1
XFILLER_200_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16193_ _08284_ _08579_ _08727_ vssd1 vssd1 vccd1 vccd1 _08838_ sky130_fd_sc_hd__o21a_1
X_15144_ _07742_ rbzero.debug_overlay.vplaneX\[-4\] vssd1 vssd1 vccd1 vccd1 _07800_
+ sky130_fd_sc_hd__nor2_1
X_12356_ net124 _05082_ _05087_ net29 net28 vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__a2111oi_2
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] _04086_ vssd1 vssd1 vccd1 vccd1
+ _04087_ sky130_fd_sc_hd__o21ai_1
X_19952_ rbzero.pov.ready_buffer\[33\] _03240_ _03243_ rbzero.debug_overlay.facingX\[-9\]
+ _03209_ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__o221a_1
X_15075_ rbzero.debug_overlay.vplaneX\[-5\] rbzero.debug_overlay.vplaneX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__or2_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12287_ net38 _05043_ _05044_ net48 vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__a22o_1
XFILLER_141_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18903_ _02558_ _02572_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__nand2_1
X_14026_ _05855_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__nand3_2
X_11238_ gpout0.hpos\[4\] vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__buf_4
X_19883_ rbzero.pov.ready_buffer\[73\] _03164_ _03155_ _03190_ vssd1 vssd1 vccd1 vccd1
+ _03191_ sky130_fd_sc_hd__o211a_1
XFILLER_150_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18834_ _02503_ _02505_ _02504_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__o21bai_1
XFILLER_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11169_ rbzero.othery\[3\] vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__inv_2
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18765_ _02450_ _02451_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__or2b_1
XFILLER_49_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15977_ _08601_ _08602_ vssd1 vssd1 vccd1 vccd1 _08622_ sky130_fd_sc_hd__xnor2_2
X_17716_ _10233_ _10280_ vssd1 vssd1 vccd1 vccd1 _10281_ sky130_fd_sc_hd__xnor2_1
X_14928_ rbzero.wall_tracer.trackDistY\[1\] rbzero.wall_tracer.trackDistX\[1\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__mux2_1
X_18696_ rbzero.wall_tracer.trackDistX\[11\] rbzero.wall_tracer.stepDistX\[11\] vssd1
+ vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__xor2_1
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17647_ _10209_ _10210_ vssd1 vssd1 vccd1 vccd1 _10212_ sky130_fd_sc_hd__and2_1
XFILLER_24_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14859_ _07576_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_21_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17578_ _10127_ _10143_ vssd1 vssd1 vccd1 vccd1 _10144_ sky130_fd_sc_hd__nand2_1
XFILLER_16_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19317_ rbzero.spi_registers.new_vshift\[1\] rbzero.spi_registers.spi_buffer\[1\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__mux2_1
XFILLER_189_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16529_ _09171_ _09172_ vssd1 vssd1 vccd1 vccd1 _09173_ sky130_fd_sc_hd__xor2_1
XFILLER_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19248_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_sky\[2\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__mux2_1
XFILLER_104_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19179_ rbzero.floor_leak\[0\] _02732_ _02734_ _02722_ vssd1 vssd1 vccd1 vccd1 _00740_
+ sky130_fd_sc_hd__o211a_1
X_21210_ clknet_leaf_30_i_clk _00979_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21141_ clknet_leaf_98_i_clk _00910_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21072_ net162 _00841_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_141_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20023_ _04992_ _04037_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__nand2_1
XFILLER_115_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20925_ clknet_leaf_74_i_clk _00694_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20856_ clknet_leaf_4_i_clk _00625_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vinf
+ sky130_fd_sc_hd__dfxtp_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20787_ clknet_leaf_47_i_clk _00556_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10540_ rbzero.tex_r0\[20\] rbzero.tex_r0\[19\] _03602_ vssd1 vssd1 vccd1 vccd1 _03607_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ rbzero.tex_r0\[53\] rbzero.tex_r0\[52\] _03569_ vssd1 vssd1 vccd1 vccd1 _03571_
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12210_ _04961_ _04960_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__and2b_1
X_21408_ net329 _01177_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13190_ _05814_ _05821_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a21oi_1
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12141_ _04909_ net62 _04911_ net12 vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__o211a_1
XFILLER_123_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21339_ net260 _01108_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[46\] sky130_fd_sc_hd__dfxtp_1
X_12072_ _04840_ _04325_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__nor2_1
XFILLER_151_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15900_ _08511_ _08543_ vssd1 vssd1 vccd1 vccd1 _08545_ sky130_fd_sc_hd__nor2_1
X_11023_ _03860_ vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__clkbuf_1
X_16880_ _08282_ _07994_ _08035_ _08046_ vssd1 vssd1 vccd1 vccd1 _09521_ sky130_fd_sc_hd__or4_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _07995_ _07989_ _08475_ vssd1 vssd1 vccd1 vccd1 _08476_ sky130_fd_sc_hd__or3_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ _02144_ _02246_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__xnor2_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _08403_ _08404_ _08405_ vssd1 vssd1 vccd1 vccd1 _08407_ sky130_fd_sc_hd__nand3_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12974_ _05586_ _05587_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__or2_2
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ _10057_ _10066_ vssd1 vssd1 vccd1 vccd1 _10067_ sky130_fd_sc_hd__nand2_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14713_ _05779_ _07362_ _07372_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__o21ai_1
X_18481_ _02176_ _02178_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__or2_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ rbzero.tex_b0\[63\] rbzero.tex_b0\[62\] _04263_ vssd1 vssd1 vccd1 vccd1 _04701_
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _07938_ _07939_ _08109_ vssd1 vssd1 vccd1 vccd1 _08338_ sky130_fd_sc_hd__or3_1
XFILLER_18_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _08747_ _09699_ _08250_ vssd1 vssd1 vccd1 vccd1 _09999_ sky130_fd_sc_hd__o21ai_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ rbzero.tex_g1\[9\] rbzero.tex_g1\[8\] _04350_ vssd1 vssd1 vccd1 vccd1 _04633_
+ sky130_fd_sc_hd__mux2_1
XFILLER_127_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14644_ _07350_ _07360_ _05793_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__mux2_1
XFILLER_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10807_ _03747_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__clkbuf_1
X_17363_ _09368_ _09217_ vssd1 vssd1 vccd1 vccd1 _09930_ sky130_fd_sc_hd__nor2_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14575_ _07305_ _07095_ _07096_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__and3_1
X_11787_ rbzero.tex_g0\[49\] rbzero.tex_g0\[48\] _04262_ vssd1 vssd1 vccd1 vccd1 _04565_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19102_ _02684_ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__clkbuf_1
X_16314_ _08290_ _08291_ _08958_ vssd1 vssd1 vccd1 vccd1 _08959_ sky130_fd_sc_hd__a21bo_1
XFILLER_174_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10738_ rbzero.tex_g0\[54\] rbzero.tex_g0\[53\] _03706_ vssd1 vssd1 vccd1 vccd1 _03711_
+ sky130_fd_sc_hd__mux2_1
X_13526_ _06256_ _06257_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__o21ai_1
X_17294_ _09854_ _09856_ _09855_ vssd1 vssd1 vccd1 vccd1 _09866_ sky130_fd_sc_hd__o21bai_1
XFILLER_203_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19033_ rbzero.pov.spi_buffer\[48\] rbzero.pov.ready_buffer\[48\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02648_ sky130_fd_sc_hd__mux2_1
X_16245_ _08881_ _08882_ vssd1 vssd1 vccd1 vccd1 _08890_ sky130_fd_sc_hd__nor2_1
X_13457_ _06152_ _06188_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__or2b_1
X_10669_ rbzero.tex_g1\[22\] rbzero.tex_g1\[23\] _03669_ vssd1 vssd1 vccd1 vccd1 _03675_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12408_ _05141_ _05172_ _05174_ net35 vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__o211a_1
XFILLER_173_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16176_ _08674_ vssd1 vssd1 vccd1 vccd1 _08821_ sky130_fd_sc_hd__clkbuf_4
X_13388_ _06046_ _06123_ _06122_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__a21bo_1
XFILLER_154_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12339_ net27 net26 vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__and2b_1
X_15127_ _07758_ _07769_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__nand2_1
XFILLER_142_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15058_ rbzero.debug_overlay.vplaneX\[-6\] _07708_ vssd1 vssd1 vccd1 vccd1 _07720_
+ sky130_fd_sc_hd__xor2_1
X_19935_ rbzero.debug_overlay.playerY\[3\] _03193_ _03229_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _01001_ sky130_fd_sc_hd__a211o_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _06240_ _06707_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__nor2_1
X_19866_ rbzero.debug_overlay.playerX\[1\] _03167_ rbzero.debug_overlay.playerX\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__o21ai_1
XFILLER_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18817_ rbzero.wall_tracer.trackDistY\[3\] rbzero.wall_tracer.stepDistY\[3\] vssd1
+ vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__nand2_1
XFILLER_56_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19599__54 clknet_1_0__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__inv_2
X_19797_ _03127_ vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18748_ _02428_ _02430_ _02429_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__a21boi_1
Xclkbuf_1_1__f__03297_ clknet_0__03297_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03297_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18679_ _02364_ _02374_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20710_ clknet_leaf_61_i_clk _00001_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.state\[3\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20641_ clknet_leaf_55_i_clk _00425_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20572_ _02721_ _03445_ _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__and3_1
XFILLER_192_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21124_ clknet_leaf_95_i_clk _00893_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21055_ clknet_leaf_1_i_clk _00824_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20006_ rbzero.pov.ready_buffer\[10\] _03239_ _03242_ _02906_ _02730_ vssd1 vssd1
+ vccd1 vccd1 _01047_ sky130_fd_sc_hd__o221a_1
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11710_ gpout0.vpos\[4\] gpout0.vpos\[3\] _04488_ gpout0.vpos\[5\] vssd1 vssd1 vccd1
+ vccd1 _04489_ sky130_fd_sc_hd__or4b_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ clknet_leaf_92_i_clk _00677_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _05435_ _05436_ _05437_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__or3b_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11641_ _04004_ _04419_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__and3b_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20839_ clknet_leaf_55_i_clk _00608_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14360_ _06882_ _07034_ _07096_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11572_ rbzero.tex_r1\[2\] _04350_ _04217_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__a21o_1
XFILLER_183_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ _06044_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__xor2_1
XFILLER_35_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10523_ rbzero.tex_r0\[28\] rbzero.tex_r0\[27\] _03591_ vssd1 vssd1 vccd1 vccd1 _03598_
+ sky130_fd_sc_hd__mux2_1
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput19 i_gpout2_sel[5] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_6
XFILLER_167_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14291_ _06798_ _06816_ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__or2b_1
XFILLER_6_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13242_ _05856_ _05877_ _05888_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__a21oi_1
X_16030_ _07980_ _08674_ _08020_ vssd1 vssd1 vccd1 vccd1 _08675_ sky130_fd_sc_hd__or3_2
XFILLER_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10454_ rbzero.tex_r0\[61\] rbzero.tex_r0\[60\] _03558_ vssd1 vssd1 vccd1 vccd1 _03562_
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13173_ _05909_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__inv_2
X_10385_ _03523_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12124_ net52 _04853_ _04857_ net50 _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__a221o_1
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17981_ _01677_ _01683_ rbzero.wall_tracer.trackDistX\[4\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00593_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19720_ _03087_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__clkbuf_1
X_16932_ _09425_ _09438_ _09572_ vssd1 vssd1 vccd1 vccd1 _09573_ sky130_fd_sc_hd__a21o_1
X_12055_ _04820_ _04823_ _04825_ _04827_ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__o32a_1
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__03320_ _03320_ vssd1 vssd1 vccd1 vccd1 clknet_0__03320_ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11006_ _03851_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19651_ _03051_ vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__clkbuf_1
X_16863_ _09502_ _09503_ vssd1 vssd1 vccd1 vccd1 _09504_ sky130_fd_sc_hd__and2b_1
XFILLER_77_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18602_ _02293_ _02298_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__xor2_1
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15814_ _08456_ _08457_ _08458_ vssd1 vssd1 vccd1 vccd1 _08459_ sky130_fd_sc_hd__a21oi_1
X_19582_ clknet_1_0__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__buf_1
X_16794_ _09428_ _09435_ vssd1 vssd1 vccd1 vccd1 _09436_ sky130_fd_sc_hd__xnor2_2
XFILLER_168_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18533_ _02132_ _02134_ _02133_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__o21bai_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _08382_ _08388_ _08389_ vssd1 vssd1 vccd1 vccd1 _08390_ sky130_fd_sc_hd__a21o_1
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _05691_ _05673_ _05683_ _05693_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__or4_2
XFILLER_46_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20060__98 clknet_1_0__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__inv_2
X_18464_ _02033_ _02055_ _02031_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a21oi_1
X_11908_ rbzero.tex_b0\[19\] rbzero.tex_b0\[18\] _04271_ vssd1 vssd1 vccd1 vccd1 _04684_
+ sky130_fd_sc_hd__mux2_1
XFILLER_206_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15676_ _08287_ _08285_ vssd1 vssd1 vccd1 vccd1 _08321_ sky130_fd_sc_hd__nand2_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12888_ rbzero.wall_tracer.visualWallDist\[2\] _05571_ _04001_ vssd1 vssd1 vccd1
+ vccd1 _05625_ sky130_fd_sc_hd__a21oi_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _09686_ _09980_ _09981_ vssd1 vssd1 vccd1 vccd1 _09982_ sky130_fd_sc_hd__a21o_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14627_ _07309_ _07310_ _07312_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__a21oi_1
X_18395_ _01859_ _01863_ _01958_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a21oi_1
X_11839_ rbzero.tex_g1\[47\] _04327_ _04328_ _04265_ vssd1 vssd1 vccd1 vccd1 _04616_
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17346_ _09633_ _09636_ _09911_ vssd1 vssd1 vccd1 vccd1 _09913_ sky130_fd_sc_hd__and3_1
XFILLER_159_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14558_ _07286_ _07292_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__xnor2_1
XFILLER_174_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13509_ _05983_ _06245_ _06243_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17277_ _05531_ _09076_ vssd1 vssd1 vccd1 vccd1 _09851_ sky130_fd_sc_hd__nand2_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14489_ _07172_ _07221_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__a21oi_1
XFILLER_146_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19016_ _02639_ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_173_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16228_ _08180_ vssd1 vssd1 vccd1 vccd1 _08873_ sky130_fd_sc_hd__clkbuf_4
XFILLER_173_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16159_ _08766_ _08800_ vssd1 vssd1 vccd1 vccd1 _08804_ sky130_fd_sc_hd__xnor2_1
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19918_ rbzero.debug_overlay.playerY\[0\] _08030_ vssd1 vssd1 vccd1 vccd1 _03216_
+ sky130_fd_sc_hd__or2_1
XFILLER_111_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19849_ _03139_ _03162_ _03163_ _03157_ vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__o211a_1
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20125__157 clknet_1_1__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__inv_2
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20624_ clknet_leaf_15_i_clk _00408_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f3 sky130_fd_sc_hd__dfxtp_2
XFILLER_178_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20555_ rbzero.traced_texVinit\[0\] _09770_ _09771_ _09068_ vssd1 vssd1 vccd1 vccd1
+ _01408_ sky130_fd_sc_hd__a22o_1
XFILLER_138_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20486_ _03383_ _03384_ _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__a21o_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21107_ net197 _00876_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21038_ clknet_leaf_75_i_clk _00807_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13860_ _06595_ _06596_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__nand2_1
X_19578__35 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__inv_2
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12811_ _05548_ _05549_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__o21bai_1
XFILLER_76_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13791_ _05824_ _06031_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__nor2_1
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15530_ _05194_ _08172_ _08174_ _08002_ vssd1 vssd1 vccd1 vccd1 _08175_ sky130_fd_sc_hd__a211o_1
XFILLER_16_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _05445_ _05489_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__xnor2_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15461_ _08086_ _08087_ _08105_ vssd1 vssd1 vccd1 vccd1 _08106_ sky130_fd_sc_hd__and3_1
X_12673_ _05419_ _05420_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__and2b_1
XFILLER_30_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17200_ rbzero.wall_tracer.mapX\[7\] _05525_ vssd1 vssd1 vccd1 vccd1 _09784_ sky130_fd_sc_hd__nor2_1
XFILLER_179_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11624_ rbzero.tex_r1\[35\] rbzero.tex_r1\[34\] _04350_ vssd1 vssd1 vccd1 vccd1 _04403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _06696_ _06698_ _07072_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__a21oi_1
X_18180_ _01879_ _01880_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__xor2_1
XFILLER_129_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15392_ _07502_ _08036_ _07933_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__mux2_4
XFILLER_169_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17131_ _03477_ _04446_ vssd1 vssd1 vccd1 vccd1 _09761_ sky130_fd_sc_hd__nand2_1
XFILLER_129_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11555_ rbzero.tex_r1\[9\] rbzero.tex_r1\[8\] _04291_ vssd1 vssd1 vccd1 vccd1 _04334_
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14343_ _07070_ _07079_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10506_ rbzero.tex_r0\[36\] rbzero.tex_r0\[35\] _03580_ vssd1 vssd1 vccd1 vccd1 _03589_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_1140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17062_ _09694_ _09701_ vssd1 vssd1 vccd1 vccd1 _09702_ sky130_fd_sc_hd__xor2_4
XFILLER_156_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14274_ _07009_ _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__xnor2_1
XFILLER_184_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11486_ _04265_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__clkbuf_8
XFILLER_100_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13225_ _05945_ _05949_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a21oi_2
X_16013_ _08656_ _08657_ vssd1 vssd1 vccd1 vccd1 _08658_ sky130_fd_sc_hd__xor2_2
XFILLER_170_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10437_ rbzero.tex_r1\[2\] rbzero.tex_r1\[3\] _03549_ vssd1 vssd1 vccd1 vccd1 _03551_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13156_ _05801_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__clkbuf_4
X_10368_ _03514_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__clkbuf_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ net3 net4 net5 vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__a21oi_1
XFILLER_135_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17964_ _01664_ _01666_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__or2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13087_ _05823_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__clkbuf_4
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10299_ _03473_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__buf_4
XFILLER_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19703_ _03078_ vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__clkbuf_1
X_12038_ _04809_ _04810_ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__o21ba_1
X_16915_ _08873_ _09555_ _09421_ vssd1 vssd1 vccd1 vccd1 _09556_ sky130_fd_sc_hd__or3b_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17895_ _01596_ _01597_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_0__03303_ _03303_ vssd1 vssd1 vccd1 vccd1 clknet_0__03303_ sky130_fd_sc_hd__clkbuf_16
XFILLER_77_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16846_ _09485_ _09486_ vssd1 vssd1 vccd1 vccd1 _09487_ sky130_fd_sc_hd__nand2_1
XFILLER_207_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19565_ rbzero.pov.spi_counter\[5\] _03031_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__and2_1
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16777_ _08237_ _09279_ _08180_ vssd1 vssd1 vccd1 vccd1 _09419_ sky130_fd_sc_hd__a21o_1
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13989_ _06725_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__inv_2
XFILLER_207_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18516_ _02109_ _02213_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__xor2_2
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15728_ _08306_ _08310_ vssd1 vssd1 vccd1 vccd1 _08373_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19496_ _02973_ _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__nand2_1
XFILLER_178_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18447_ _01737_ _10238_ _09292_ _09991_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__or4_1
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15659_ _08255_ _08303_ vssd1 vssd1 vccd1 vccd1 _08304_ sky130_fd_sc_hd__nand2_1
XFILLER_178_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18378_ _01474_ _09215_ _01941_ _02076_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__o31a_1
XFILLER_159_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17329_ _09896_ vssd1 vssd1 vccd1 vccd1 _09897_ sky130_fd_sc_hd__inv_2
XFILLER_105_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20271_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__buf_1
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21656_ clknet_leaf_90_i_clk _01425_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20607_ gpout3.clk_div\[1\] gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__or2_1
XFILLER_162_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21587_ net508 _01356_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_75 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_75/HI o_rgb[3] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_86 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_86/HI o_rgb[18] sky130_fd_sc_hd__conb_1
XFILLER_165_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ _04099_ _04069_ _04097_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__nor3_2
Xtop_ew_algofoogle_97 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_97/HI zeros[7] sky130_fd_sc_hd__conb_1
X_20538_ rbzero.texV\[8\] _03327_ _03332_ _03429_ vssd1 vssd1 vccd1 vccd1 _01404_
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11271_ _04049_ _04050_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__nand2_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20469_ _03272_ _03370_ _03371_ _03250_ rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1
+ _01393_ sky130_fd_sc_hd__a32o_1
X_13010_ _05690_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__inv_2
XFILLER_134_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14961_ _05201_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__buf_4
XFILLER_181_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16700_ _09324_ _09326_ vssd1 vssd1 vccd1 vccd1 _09342_ sky130_fd_sc_hd__or2_2
XFILLER_43_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13912_ _06576_ _06648_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__nand2_1
XFILLER_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17680_ _10099_ _10244_ vssd1 vssd1 vccd1 vccd1 _10245_ sky130_fd_sc_hd__xnor2_2
XFILLER_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14892_ _07602_ _04019_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__nand2_1
XFILLER_63_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16631_ _09269_ _09273_ vssd1 vssd1 vccd1 vccd1 _09274_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13843_ _06259_ _06575_ _06578_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__or3_1
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19350_ rbzero.debug_overlay.vplaneY\[-4\] rbzero.wall_tracer.rayAddendY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__nor2_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20108__141 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__inv_2
X_16562_ _09059_ _08470_ _08546_ vssd1 vssd1 vccd1 vccd1 _09205_ sky130_fd_sc_hd__or3_1
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10986_ net48 rbzero.tex_b0\[63\] _03762_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__mux2_1
X_13774_ _05944_ _06009_ _06510_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__or3b_1
X_18301_ _01966_ _02000_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__xnor2_2
XFILLER_203_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15513_ _05208_ _08157_ vssd1 vssd1 vccd1 vccd1 _08158_ sky130_fd_sc_hd__or2_1
XFILLER_204_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12725_ _05424_ _05425_ _05427_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__o21a_1
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19281_ _02795_ vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16493_ _08981_ _07574_ _08234_ _09136_ _07970_ vssd1 vssd1 vccd1 vccd1 _09137_ sky130_fd_sc_hd__a311o_1
XFILLER_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18232_ _01930_ _01931_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__nand2_1
XFILLER_31_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15444_ _08030_ _08088_ vssd1 vssd1 vccd1 vccd1 _08089_ sky130_fd_sc_hd__and2_1
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12656_ _05388_ _05398_ _05399_ _05397_ rbzero.map_rom.i_row\[4\] vssd1 vssd1 vccd1
+ vccd1 _05406_ sky130_fd_sc_hd__a32o_1
XFILLER_141_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18163_ _01739_ _01620_ _01862_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__o21ai_1
X_11607_ _04384_ _04385_ _04226_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__mux2_1
X_12587_ _05323_ _05288_ _05319_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__or3_1
X_15375_ _05197_ rbzero.wall_tracer.stepDistX\[-7\] vssd1 vssd1 vccd1 vccd1 _08020_
+ sky130_fd_sc_hd__nor2_1
XFILLER_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17114_ _04821_ _09750_ _09751_ vssd1 vssd1 vccd1 vccd1 _09752_ sky130_fd_sc_hd__and3_1
X_14326_ _06240_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__and3b_1
X_11538_ _04317_ _04163_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__and2_1
X_18094_ _01793_ _01794_ _01795_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__a21oi_1
XFILLER_184_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17045_ _09141_ _09420_ _08194_ vssd1 vssd1 vccd1 vccd1 _09685_ sky130_fd_sc_hd__a21o_1
X_11469_ rbzero.tex_r0\[43\] rbzero.tex_r0\[42\] _04213_ vssd1 vssd1 vccd1 vccd1 _04249_
+ sky130_fd_sc_hd__mux2_1
X_14257_ _06884_ _06915_ _06917_ _06993_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__or4_2
XFILLER_7_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20154__183 clknet_1_0__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__inv_2
X_13208_ _05856_ _05877_ _05944_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__a21o_2
X_14188_ _06769_ _06671_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__nor2_1
XFILLER_140_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ _05865_ _05870_ _05875_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__or3b_1
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ rbzero.pov.spi_buffer\[30\] rbzero.pov.ready_buffer\[30\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02629_ sky130_fd_sc_hd__mux2_1
XFILLER_112_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _01647_ _01648_ _01649_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__and3_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17878_ _09661_ _09029_ _09165_ _01462_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__o22ai_1
XFILLER_66_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16829_ _09461_ _09465_ vssd1 vssd1 vccd1 vccd1 _09470_ sky130_fd_sc_hd__or2_1
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19548_ rbzero.pov.spi_counter\[0\] _03019_ _03021_ vssd1 vssd1 vccd1 vccd1 _00822_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_94_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19479_ _02941_ _02944_ _02957_ _02959_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__o31a_1
XFILLER_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21510_ net431 _01279_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21441_ net362 _01210_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20237__258 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__inv_2
XFILLER_119_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21372_ net293 _01141_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_i_clk clknet_3_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10840_ rbzero.tex_g0\[6\] rbzero.tex_g0\[5\] _03762_ vssd1 vssd1 vccd1 vccd1 _03765_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ _03728_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ rbzero.wall_tracer.trackDistY\[3\] _05264_ rbzero.wall_tracer.trackDistY\[-5\]
+ _05236_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a22o_1
X_13490_ _06225_ _06226_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__and2_1
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ net71 rbzero.wall_tracer.state\[5\] _05190_ vssd1 vssd1 vccd1 vccd1 _05199_
+ sky130_fd_sc_hd__and3_1
XFILLER_12_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21639_ clknet_leaf_28_i_clk _01408_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12372_ net33 net32 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__nor2_2
X_15160_ _07803_ _07808_ _07813_ _07676_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__o31ai_1
Xclkbuf_leaf_43_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_197_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11323_ rbzero.texV\[8\] _04102_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__xor2_1
X_14111_ _06843_ _06844_ _06846_ _06847_ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__a22o_1
XFILLER_153_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15091_ _07736_ _07748_ _07749_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__or3_1
XFILLER_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14042_ _06002_ _06758_ _06759_ _06770_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__a31o_1
X_11254_ _04031_ _04032_ _04002_ _04035_ _00000_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__a41o_1
XFILLER_153_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18850_ _02517_ _02519_ _02518_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__o21bai_1
Xclkbuf_leaf_58_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_192_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11185_ rbzero.map_rom.f2 _03933_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__nand2_1
XFILLER_192_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17801_ _10244_ _01503_ _01504_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__a21o_1
XFILLER_67_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18781_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__and2_1
X_15993_ _08629_ _08637_ vssd1 vssd1 vccd1 vccd1 _08638_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17732_ _10295_ _10296_ vssd1 vssd1 vccd1 vccd1 _10297_ sky130_fd_sc_hd__and2b_2
XFILLER_76_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14944_ rbzero.wall_tracer.visualWallDist\[6\] _07618_ vssd1 vssd1 vccd1 vccd1 _07639_
+ sky130_fd_sc_hd__or2_1
XFILLER_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17663_ _10225_ _10227_ vssd1 vssd1 vccd1 vccd1 _10228_ sky130_fd_sc_hd__nor2_1
X_14875_ _05737_ _05736_ _07588_ _07468_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__nor4_4
XFILLER_169_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19402_ _02886_ _02887_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__and2_1
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16614_ _09009_ _09099_ vssd1 vssd1 vccd1 vccd1 _09257_ sky130_fd_sc_hd__nand2_1
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13826_ _06335_ _06560_ _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__a21oi_4
X_17594_ _10048_ _10159_ vssd1 vssd1 vccd1 vccd1 _10160_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19333_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.wall_tracer.rayAddendY\[-5\] vssd1
+ vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__nor2_1
X_16545_ _09055_ vssd1 vssd1 vccd1 vccd1 _09189_ sky130_fd_sc_hd__inv_2
X_13757_ _06438_ _06455_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__xor2_1
XFILLER_91_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10969_ _03832_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12708_ _05447_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__xor2_4
X_19264_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_floor\[2\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__mux2_1
XFILLER_206_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16476_ _08283_ _08177_ _08264_ _08626_ vssd1 vssd1 vccd1 vccd1 _09120_ sky130_fd_sc_hd__a2bb2o_1
X_13688_ _06376_ _06424_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__or2b_1
X_18215_ _01897_ _01899_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__or2_1
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15427_ _07904_ _08071_ vssd1 vssd1 vccd1 vccd1 _08072_ sky130_fd_sc_hd__nand2_1
X_19195_ _09753_ _02743_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__and2_1
X_12639_ _05388_ _05390_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__nand2_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18146_ _01840_ _01846_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__xnor2_2
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15358_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\] rbzero.debug_overlay.playerY\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _08003_ sky130_fd_sc_hd__o21ai_1
XFILLER_172_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14309_ _06696_ _06667_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__nor2_1
X_18077_ _01611_ _01655_ _01778_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__a21oi_1
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15289_ _05349_ _05469_ rbzero.wall_tracer.side vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__mux2_1
XFILLER_89_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17028_ _08570_ vssd1 vssd1 vccd1 vccd1 _09668_ sky130_fd_sc_hd__buf_4
XFILLER_132_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18979_ rbzero.pov.spi_buffer\[22\] rbzero.pov.ready_buffer\[22\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02620_ sky130_fd_sc_hd__mux2_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20941_ clknet_leaf_3_i_clk _00710_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_54_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20872_ clknet_leaf_95_i_clk _00641_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21424_ net345 _01193_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21355_ net276 _01124_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21286_ clknet_leaf_36_i_clk _01055_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[4\] sky130_fd_sc_hd__dfxtp_4
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _05724_ _05683_ _05726_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__o21ba_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11941_ rbzero.tex_b0\[43\] rbzero.tex_b0\[42\] _04342_ vssd1 vssd1 vccd1 vccd1 _04717_
+ sky130_fd_sc_hd__mux2_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _07371_ _07396_ _05779_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__mux2_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ rbzero.tex_g1\[21\] rbzero.tex_g1\[20\] _04336_ vssd1 vssd1 vccd1 vccd1 _04649_
+ sky130_fd_sc_hd__mux2_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _06304_ _06323_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__xnor2_1
X_10823_ rbzero.tex_g0\[14\] rbzero.tex_g0\[13\] _03751_ vssd1 vssd1 vccd1 vccd1 _03756_
+ sky130_fd_sc_hd__mux2_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14591_ _07326_ _07327_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__xnor2_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ _08178_ _08194_ vssd1 vssd1 vccd1 vccd1 _08975_ sky130_fd_sc_hd__nor2_1
XFILLER_129_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13542_ _06150_ _06192_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__xnor2_2
XFILLER_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10754_ rbzero.tex_g0\[47\] rbzero.tex_g0\[46\] _03718_ vssd1 vssd1 vccd1 vccd1 _03720_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _08902_ _08904_ vssd1 vssd1 vccd1 vccd1 _08906_ sky130_fd_sc_hd__nand2_1
X_10685_ _03683_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__clkbuf_1
X_13473_ _06165_ _06158_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__or2b_1
XFILLER_200_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18000_ _09526_ _01576_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__nor2_1
XFILLER_185_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15212_ _07820_ rbzero.wall_tracer.rayAddendX\[8\] vssd1 vssd1 vccd1 vccd1 _07864_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12424_ _05188_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__clkbuf_4
X_16192_ _08828_ _08829_ _08831_ vssd1 vssd1 vccd1 vccd1 _08837_ sky130_fd_sc_hd__or3b_1
XFILLER_127_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20372__379 clknet_1_0__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__inv_2
X_15143_ _07797_ _07798_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__xnor2_1
X_12355_ _05117_ _05119_ _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__and3_1
XFILLER_114_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ rbzero.traced_texVinit\[2\] rbzero.texV\[2\] rbzero.texV\[1\] rbzero.traced_texVinit\[1\]
+ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__a221o_1
X_12286_ net23 vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__inv_2
X_15074_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.debug_overlay.vplaneX\[-8\] rbzero.debug_overlay.vplaneX\[-9\]
+ rbzero.debug_overlay.vplaneX\[-5\] vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__or4b_1
X_19951_ _03242_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__buf_2
XFILLER_114_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11237_ _04020_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__buf_6
X_18902_ _02559_ rbzero.spi_registers.spi_counter\[0\] _02566_ _02568_ _02571_ vssd1
+ vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__o2111a_1
X_14025_ _06704_ _06760_ _06761_ _05825_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__o22ai_2
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19882_ _03188_ _03185_ _02822_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__a21o_1
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18833_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.stepDistY\[5\] vssd1
+ vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__nand2_1
X_11168_ rbzero.otherx\[0\] _03919_ _03935_ rbzero.othery\[4\] _03956_ vssd1 vssd1
+ vccd1 vccd1 _03957_ sky130_fd_sc_hd__a221o_1
XFILLER_110_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18764_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.stepDistY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__nand2_1
X_11099_ _03900_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__clkbuf_1
X_15976_ _08605_ _08606_ vssd1 vssd1 vccd1 vccd1 _08621_ sky130_fd_sc_hd__xnor2_2
XFILLER_82_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17715_ _10277_ _10279_ vssd1 vssd1 vccd1 vccd1 _10280_ sky130_fd_sc_hd__xnor2_1
X_20266__284 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__inv_2
XFILLER_76_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14927_ _07621_ _07626_ _07627_ _07620_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__o211a_1
X_18695_ _02319_ _02320_ _02318_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__o21ai_1
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17646_ _10209_ _10210_ vssd1 vssd1 vccd1 vccd1 _10211_ sky130_fd_sc_hd__nor2_1
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14858_ rbzero.wall_tracer.stepDistY\[7\] _07575_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07576_ sky130_fd_sc_hd__mux2_1
XFILLER_91_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13809_ _06500_ _06493_ _06544_ _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__or4b_1
X_17577_ _10140_ _10141_ _10137_ vssd1 vssd1 vccd1 vccd1 _10143_ sky130_fd_sc_hd__a21o_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14789_ _05800_ _07520_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__nand2_1
XFILLER_189_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19316_ _02814_ vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_91_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16528_ _08054_ _08425_ vssd1 vssd1 vccd1 vccd1 _09172_ sky130_fd_sc_hd__nor2_1
XFILLER_176_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19247_ _02776_ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__clkbuf_1
X_16459_ _08097_ vssd1 vssd1 vccd1 vccd1 _09103_ sky130_fd_sc_hd__clkbuf_4
XFILLER_192_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19178_ rbzero.spi_registers.new_leak\[0\] _02733_ vssd1 vssd1 vccd1 vccd1 _02734_
+ sky130_fd_sc_hd__or2_1
XFILLER_117_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18129_ _07974_ _09217_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__or2_1
XFILLER_172_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21140_ clknet_leaf_98_i_clk _00909_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21071_ net161 _00840_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_101_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20022_ _04021_ _04026_ _03266_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__and3_1
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20924_ clknet_leaf_26_i_clk _00693_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20855_ clknet_leaf_51_i_clk _00624_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20786_ clknet_leaf_47_i_clk _00555_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_179_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10470_ _03570_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21407_ net328 _01176_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12140_ _04910_ net61 vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__or2_1
XFILLER_123_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21338_ net259 _01107_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ net6 _04841_ _04842_ net5 vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a31o_1
XFILLER_173_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21269_ clknet_leaf_89_i_clk _01038_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ rbzero.tex_b0\[47\] rbzero.tex_b0\[46\] _03854_ vssd1 vssd1 vccd1 vccd1 _03860_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _07980_ _07929_ _07930_ vssd1 vssd1 vccd1 vccd1 _08475_ sky130_fd_sc_hd__or3_2
XFILLER_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _08403_ _08404_ _08405_ vssd1 vssd1 vccd1 vccd1 _08406_ sky130_fd_sc_hd__a21o_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ _05582_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__xor2_4
XFILLER_58_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17500_ _10064_ _10065_ vssd1 vssd1 vccd1 vccd1 _10066_ sky130_fd_sc_hd__and2_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _05963_ _07445_ _07446_ _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__o31a_1
XFILLER_205_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18480_ _10094_ _09215_ _02072_ _02177_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__o31a_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _04140_ _04683_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__or3_1
XFILLER_206_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15692_ _08334_ _08336_ vssd1 vssd1 vccd1 vccd1 _08337_ sky130_fd_sc_hd__xnor2_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17431_ _08377_ _08519_ _09699_ vssd1 vssd1 vccd1 vccd1 _09998_ sky130_fd_sc_hd__a21o_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _07378_ _07335_ _07336_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__or3b_1
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _04629_ _04630_ _04631_ _04379_ _04209_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__o221a_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17362_ _09927_ _09928_ vssd1 vssd1 vccd1 vccd1 _09929_ sky130_fd_sc_hd__nand2_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10806_ rbzero.tex_g0\[22\] rbzero.tex_g0\[21\] _03740_ vssd1 vssd1 vccd1 vccd1 _03747_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14574_ _07309_ _07310_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__nand2_1
XFILLER_207_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11786_ _04306_ _04559_ _04563_ _04371_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__a211o_1
XFILLER_14_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19101_ rbzero.spi_registers.spi_buffer\[6\] rbzero.spi_registers.spi_buffer\[5\]
+ _02677_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__mux2_1
XFILLER_198_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16313_ _08292_ _07996_ _07959_ vssd1 vssd1 vccd1 vccd1 _08958_ sky130_fd_sc_hd__or3_1
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13525_ _06258_ _06261_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__xnor2_1
X_10737_ _03710_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__clkbuf_1
X_17293_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.stepDistX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _09865_ sky130_fd_sc_hd__nand2_1
XFILLER_202_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19032_ _02647_ vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__clkbuf_1
X_16244_ _08827_ _08833_ vssd1 vssd1 vccd1 vccd1 _08889_ sky130_fd_sc_hd__xnor2_1
XFILLER_139_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13456_ _06150_ _06192_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__and2b_1
XFILLER_174_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ _03674_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12407_ _05145_ _05173_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__or2_1
X_16175_ _08818_ _08819_ vssd1 vssd1 vccd1 vccd1 _08820_ sky130_fd_sc_hd__or2_1
X_10599_ rbzero.tex_g1\[55\] rbzero.tex_g1\[56\] _03635_ vssd1 vssd1 vccd1 vccd1 _03638_
+ sky130_fd_sc_hd__mux2_1
X_13387_ _06122_ _06046_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__nand3b_1
XFILLER_103_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15126_ _07761_ _07771_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__nor2_1
X_12338_ net48 net39 net38 net40 _05082_ _05087_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__mux4_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15057_ _07719_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__clkbuf_1
X_19934_ rbzero.pov.ready_buffer\[56\] _03146_ _03227_ _03228_ _03197_ vssd1 vssd1
+ vccd1 vccd1 _03229_ sky130_fd_sc_hd__o221a_1
XFILLER_114_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12269_ _04989_ _04990_ _05021_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__mux2_1
XFILLER_141_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14008_ _06245_ _06668_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__nor2_1
XFILLER_96_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19865_ rbzero.debug_overlay.playerX\[2\] rbzero.debug_overlay.playerX\[1\] _03167_
+ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__or3_1
XFILLER_110_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18816_ _02496_ _01438_ rbzero.wall_tracer.trackDistY\[2\] _02406_ vssd1 vssd1 vccd1
+ vccd1 _00615_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19796_ rbzero.pov.spi_buffer\[71\] rbzero.pov.spi_buffer\[72\] _03047_ vssd1 vssd1
+ vccd1 vccd1 _03127_ sky130_fd_sc_hd__mux2_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18747_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.stepDistY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__and2_1
X_15959_ _08601_ _08602_ _08603_ vssd1 vssd1 vccd1 vccd1 _08604_ sky130_fd_sc_hd__a21oi_2
XFILLER_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03296_ clknet_0__03296_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03296_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18678_ _02367_ _02373_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17629_ _10192_ _10193_ vssd1 vssd1 vccd1 vccd1 _10194_ sky130_fd_sc_hd__nor2_1
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20640_ clknet_leaf_64_i_clk _00424_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_177_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20571_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__or2_1
XFILLER_192_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21123_ net213 _00892_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_120_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21054_ clknet_leaf_1_i_clk _00823_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20005_ rbzero.pov.ready_buffer\[9\] _03239_ _03242_ rbzero.debug_overlay.vplaneY\[0\]
+ _02730_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__o221a_1
XFILLER_87_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20907_ clknet_leaf_91_i_clk _00676_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _04022_ _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__and2b_1
XFILLER_39_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20838_ clknet_leaf_54_i_clk _00607_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_70_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20102__136 clknet_1_1__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__inv_2
XFILLER_51_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ _04336_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__clkbuf_8
X_20769_ clknet_leaf_43_i_clk _00538_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13310_ _05995_ _05921_ _06046_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__o21ai_1
XFILLER_7_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10522_ _03597_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_161_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14290_ _07006_ _07026_ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__xnor2_2
XFILLER_11_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10453_ _03561_ vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13241_ _05939_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__buf_2
XFILLER_202_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10384_ rbzero.tex_r1\[27\] rbzero.tex_r1\[28\] _03516_ vssd1 vssd1 vccd1 vccd1 _03523_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13172_ _05871_ _05905_ _05907_ _05908_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__o211a_2
XFILLER_124_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12123_ net49 _04838_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__and2_1
XFILLER_11_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17980_ _01681_ _01682_ _09780_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16931_ _09436_ _09437_ vssd1 vssd1 vccd1 vccd1 _09572_ sky130_fd_sc_hd__and2b_1
X_12054_ _03473_ rbzero.row_render.wall\[0\] _04814_ vssd1 vssd1 vccd1 vccd1 _04828_
+ sky130_fd_sc_hd__and3b_1
XFILLER_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11005_ rbzero.tex_b0\[55\] rbzero.tex_b0\[54\] _03843_ vssd1 vssd1 vccd1 vccd1 _03851_
+ sky130_fd_sc_hd__mux2_1
XFILLER_172_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16862_ _09245_ _08075_ _08159_ _08150_ vssd1 vssd1 vccd1 vccd1 _09503_ sky130_fd_sc_hd__or4_1
X_19650_ rbzero.pov.spi_buffer\[1\] rbzero.pov.spi_buffer\[2\] _03048_ vssd1 vssd1
+ vccd1 vccd1 _03051_ sky130_fd_sc_hd__mux2_1
XFILLER_77_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18601_ _02296_ _02297_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__nor2_1
X_15813_ _08442_ _08455_ vssd1 vssd1 vccd1 vccd1 _08458_ sky130_fd_sc_hd__nor2_1
X_16793_ _08239_ _09434_ vssd1 vssd1 vccd1 vccd1 _09435_ sky130_fd_sc_hd__nor2_1
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18532_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.stepDistX\[9\] vssd1
+ vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__nand2_1
XFILLER_93_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15744_ _08375_ _08381_ vssd1 vssd1 vccd1 vccd1 _08389_ sky130_fd_sc_hd__nor2_1
XFILLER_206_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12956_ _05692_ _05636_ _05648_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__or3b_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _02141_ _02160_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__xnor2_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _04232_ _04670_ _04674_ _04682_ _04244_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__o311a_1
X_15675_ _08318_ _08309_ _08319_ vssd1 vssd1 vccd1 vccd1 _08320_ sky130_fd_sc_hd__a21o_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _05333_ _05334_ _04031_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__o21ai_1
XFILLER_61_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _08767_ _09552_ _09973_ _08283_ vssd1 vssd1 vccd1 vccd1 _09981_ sky130_fd_sc_hd__o22a_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _07095_ _07035_ _07099_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__a21oi_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ _02084_ _02092_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__xnor2_1
X_11838_ rbzero.tex_g1\[46\] _04272_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__and2_1
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _09633_ _09636_ _09911_ vssd1 vssd1 vccd1 vccd1 _09912_ sky130_fd_sc_hd__a21oi_2
X_20378__385 clknet_1_1__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__inv_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _07285_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__xor2_1
XFILLER_92_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11769_ rbzero.tex_g0\[27\] rbzero.tex_g0\[26\] _04341_ vssd1 vssd1 vccd1 vccd1 _04547_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20077__113 clknet_1_1__leaf__03290_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__inv_2
XFILLER_146_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ _05940_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__clkbuf_4
XFILLER_158_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17276_ _09846_ _09847_ _09848_ vssd1 vssd1 vccd1 vccd1 _09850_ sky130_fd_sc_hd__a21oi_1
XFILLER_147_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14488_ _07222_ _07224_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__and2b_1
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19015_ rbzero.pov.spi_buffer\[39\] rbzero.pov.ready_buffer\[39\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02639_ sky130_fd_sc_hd__mux2_1
X_16227_ _08170_ vssd1 vssd1 vccd1 vccd1 _08872_ sky130_fd_sc_hd__clkbuf_4
X_13439_ _06080_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__clkinv_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16158_ _08802_ _08579_ _08777_ vssd1 vssd1 vccd1 vccd1 _08803_ sky130_fd_sc_hd__or3_1
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15109_ rbzero.wall_tracer.rayAddendX\[1\] _07695_ _07767_ _07703_ vssd1 vssd1 vccd1
+ vccd1 _07768_ sky130_fd_sc_hd__a22o_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16089_ _08726_ _08733_ vssd1 vssd1 vccd1 vccd1 _08734_ sky130_fd_sc_hd__or2b_1
XFILLER_170_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19917_ rbzero.debug_overlay.playerY\[-1\] _03193_ _03215_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _00997_ sky130_fd_sc_hd__a211o_1
XFILLER_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19848_ _08078_ _03143_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__nand2_1
XFILLER_95_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19779_ _03118_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__clkbuf_1
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20623_ clknet_leaf_15_i_clk _00407_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.f4 sky130_fd_sc_hd__dfxtp_2
XFILLER_165_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20554_ _03441_ _03442_ rbzero.texV\[11\] net60 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_192_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20485_ _03379_ _03381_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__nand2_1
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21106_ net196 _00875_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21037_ clknet_leaf_77_i_clk _00806_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ rbzero.wall_tracer.mapY\[8\] _05404_ _05547_ vssd1 vssd1 vccd1 vccd1 _05550_
+ sky130_fd_sc_hd__a21bo_1
X_13790_ _06382_ _06002_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__nand2_1
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _05416_ _05442_ _05443_ _05444_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__a31o_1
XFILLER_76_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15460_ _08097_ _08104_ vssd1 vssd1 vccd1 vccd1 _08105_ sky130_fd_sc_hd__nor2_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__nand2_1
XFILLER_70_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _07115_ _07119_ _07117_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__o21ba_1
XFILLER_187_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11623_ _04379_ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__or2_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15391_ _05355_ _05477_ _07893_ vssd1 vssd1 vccd1 vccd1 _08036_ sky130_fd_sc_hd__mux2_1
XFILLER_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17130_ _03477_ _04446_ vssd1 vssd1 vccd1 vccd1 _09760_ sky130_fd_sc_hd__or2_1
X_14342_ _07077_ _07078_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__xor2_1
XFILLER_155_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11554_ _04326_ _04330_ _04331_ _04247_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__o221a_1
XFILLER_195_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10505_ _03588_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__clkbuf_1
X_17061_ _09696_ _09700_ vssd1 vssd1 vccd1 vccd1 _09701_ sky130_fd_sc_hd__xnor2_2
XFILLER_156_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14273_ _06680_ _06708_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__nor2_1
XFILLER_13_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11485_ _04126_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__buf_6
XFILLER_143_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03299_ clknet_0__03299_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03299_
+ sky130_fd_sc_hd__clkbuf_16
X_16012_ _08578_ _08580_ vssd1 vssd1 vccd1 vccd1 _08657_ sky130_fd_sc_hd__xnor2_2
XFILLER_13_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13224_ _05800_ _05950_ _05955_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__o211a_2
XFILLER_155_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10436_ _03550_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13155_ _05743_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__clkbuf_4
X_10367_ rbzero.tex_r1\[35\] rbzero.tex_r1\[36\] _03505_ vssd1 vssd1 vccd1 vccd1 _03514_
+ sky130_fd_sc_hd__mux2_1
XFILLER_152_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _04154_ _03477_ _04840_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__mux2_1
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17963_ _01543_ _01545_ _01665_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__o21a_1
X_10298_ gpout0.hpos\[0\] vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__buf_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _05800_ _05812_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__o21ai_4
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19702_ rbzero.pov.spi_buffer\[26\] rbzero.pov.spi_buffer\[27\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03078_ sky130_fd_sc_hd__mux2_1
X_12037_ _04004_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__buf_2
X_16914_ _09554_ _09138_ _05198_ vssd1 vssd1 vccd1 vccd1 _09555_ sky130_fd_sc_hd__mux2_2
XFILLER_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17894_ _08275_ _08427_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0__03302_ _03302_ vssd1 vssd1 vccd1 vccd1 clknet_0__03302_ sky130_fd_sc_hd__clkbuf_16
X_16845_ _08160_ _09352_ _09484_ vssd1 vssd1 vccd1 vccd1 _09486_ sky130_fd_sc_hd__or3_1
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16776_ _09117_ _09417_ vssd1 vssd1 vccd1 vccd1 _09418_ sky130_fd_sc_hd__nor2_1
X_19564_ _03033_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_92_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13988_ _06696_ _06677_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__nor2_1
XFILLER_94_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18515_ _02211_ _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__nor2_1
X_15727_ _08313_ _08324_ vssd1 vssd1 vccd1 vccd1 _08372_ sky130_fd_sc_hd__xnor2_1
XFILLER_207_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12939_ _05601_ _05604_ _05638_ _05649_ _05628_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__o41a_1
XFILLER_207_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _02904_ rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 _02974_
+ sky130_fd_sc_hd__or2_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18446_ _01971_ _02027_ _02036_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__o21ai_4
X_15658_ rbzero.wall_tracer.visualWallDist\[-11\] _08148_ _05198_ _08199_ vssd1 vssd1
+ vccd1 vccd1 _08303_ sky130_fd_sc_hd__and4_1
XFILLER_179_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14609_ _07218_ _07323_ _07334_ _07332_ _07345_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__a311o_1
X_18377_ _01939_ _01940_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__nand2_1
XFILLER_159_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15589_ _08218_ _08232_ _08208_ vssd1 vssd1 vccd1 vccd1 _08234_ sky130_fd_sc_hd__and3_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17328_ _04016_ _09739_ vssd1 vssd1 vccd1 vccd1 _09896_ sky130_fd_sc_hd__nand2_1
XFILLER_146_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17259_ _05531_ _09069_ vssd1 vssd1 vccd1 vccd1 _09835_ sky130_fd_sc_hd__nand2_1
XFILLER_190_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20131__162 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__inv_2
XFILLER_64_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21655_ clknet_leaf_90_i_clk _01424_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20606_ gpout3.clk_div\[1\] gpout3.clk_div\[0\] vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__nand2_1
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21586_ net507 _01355_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_193_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_76 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_76/HI o_rgb[4] sky130_fd_sc_hd__conb_1
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xtop_ew_algofoogle_87 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_87/HI o_rgb[19] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_98 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_98/HI zeros[8] sky130_fd_sc_hd__conb_1
X_20537_ _03426_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11270_ rbzero.traced_texVinit\[10\] rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1 _04050_
+ sky130_fd_sc_hd__or2_1
X_20468_ _03367_ _03368_ _03369_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nand3_1
XFILLER_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20214__237 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__inv_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14960_ rbzero.wall_tracer.visualWallDist\[11\] _07595_ _07649_ _07642_ vssd1 vssd1
+ vccd1 vccd1 _00466_ sky130_fd_sc_hd__o211a_1
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13911_ _06569_ _06647_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__xnor2_1
XFILLER_101_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14891_ _07601_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__clkinv_2
XFILLER_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16630_ _09271_ _09272_ vssd1 vssd1 vccd1 vccd1 _09273_ sky130_fd_sc_hd__xnor2_1
X_13842_ _06259_ _06575_ _06578_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16561_ _09059_ _09193_ vssd1 vssd1 vccd1 vccd1 _09204_ sky130_fd_sc_hd__and2b_1
X_13773_ _05823_ _06045_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__nor2_1
X_10985_ _03840_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18300_ _01998_ _01999_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__xor2_2
XFILLER_71_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15512_ rbzero.wall_tracer.visualWallDist\[4\] _08148_ vssd1 vssd1 vccd1 vccd1 _08157_
+ sky130_fd_sc_hd__nand2_4
X_12724_ _05470_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__xnor2_2
X_19280_ rbzero.spi_registers.spi_buffer\[2\] rbzero.spi_registers.new_leak\[2\] _02792_
+ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__mux2_1
XFILLER_204_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16492_ _07566_ _07568_ _07571_ _08220_ _07575_ vssd1 vssd1 vccd1 vccd1 _09136_ sky130_fd_sc_hd__o41a_1
XFILLER_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20295__309 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__inv_2
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18231_ _01875_ _01857_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__or2b_1
XFILLER_188_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15443_ rbzero.debug_overlay.playerY\[-2\] _08029_ rbzero.debug_overlay.playerY\[-1\]
+ vssd1 vssd1 vccd1 vccd1 _08088_ sky130_fd_sc_hd__o21ai_1
X_12655_ rbzero.wall_tracer.mapY\[5\] _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__xnor2_1
XFILLER_90_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18162_ _01739_ _01620_ _01862_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__or3_1
X_11606_ rbzero.tex_r1\[51\] rbzero.tex_r1\[50\] _04338_ vssd1 vssd1 vccd1 vccd1 _04385_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15374_ _04013_ _08017_ _08018_ vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__a21oi_2
XFILLER_90_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12586_ _05338_ _05339_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__and2_1
XFILLER_8_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17113_ _04814_ _03474_ vssd1 vssd1 vccd1 vccd1 _09751_ sky130_fd_sc_hd__or2_1
X_14325_ _06245_ _06708_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__or2_1
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11537_ gpout0.hpos\[2\] vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__clkbuf_4
X_18093_ _01678_ _01680_ _01679_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__o21bai_1
XFILLER_8_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17044_ _08767_ _09417_ vssd1 vssd1 vccd1 vccd1 _09684_ sky130_fd_sc_hd__nor2_1
XFILLER_172_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14256_ _06982_ _06989_ _06991_ _06992_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__a211oi_1
XFILLER_183_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11468_ _04245_ _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__mux2_1
XFILLER_172_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13207_ _05700_ _05879_ _05881_ _05887_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__a211o_1
X_10419_ _03541_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__clkbuf_1
X_14187_ _06894_ _06896_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__xnor2_1
XFILLER_87_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11399_ _04153_ _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__nor2_1
X_20189__214 clknet_1_0__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__inv_2
XFILLER_135_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _05703_ _05871_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__or3_1
XFILLER_140_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _02628_ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17946_ _01523_ _01529_ _10271_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__a21o_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _05777_ _05796_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__xnor2_1
XFILLER_79_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17877_ _01578_ _01579_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__xnor2_1
XFILLER_65_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16828_ rbzero.wall_tracer.texu\[3\] _09085_ _09468_ _09469_ _07642_ vssd1 vssd1
+ vccd1 vccd1 _00514_ sky130_fd_sc_hd__o221a_1
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19547_ rbzero.pov.spi_counter\[0\] _03019_ _03020_ vssd1 vssd1 vccd1 vccd1 _03021_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_111_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16759_ _09252_ _09394_ _09399_ vssd1 vssd1 vccd1 vccd1 _09401_ sky130_fd_sc_hd__and3_1
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19478_ _04034_ _02958_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__nor2_1
XFILLER_55_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18429_ _01799_ _02024_ _02025_ _02023_ _02127_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__a221o_4
XFILLER_142_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21440_ net361 _01209_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21371_ net292 _01140_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19635__87 clknet_1_0__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__inv_2
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10770_ rbzero.tex_g0\[39\] rbzero.tex_g0\[38\] _03718_ vssd1 vssd1 vccd1 vccd1 _03728_
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_922 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12440_ _05198_ _03914_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__nor2_1
XFILLER_185_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21638_ clknet_leaf_40_i_clk _01407_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12371_ net35 net36 net37 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__nor3_2
XFILLER_165_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21569_ net490 _01338_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14110_ _06666_ _06678_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__nor2_1
XFILLER_138_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11322_ _04055_ _04054_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__nand2_1
X_15090_ _07748_ _07749_ _07736_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__o21ai_1
XFILLER_165_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14041_ _06012_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__and3_1
XFILLER_107_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11253_ _04034_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__buf_4
X_11184_ rbzero.map_rom.f2 rbzero.map_rom.f1 rbzero.map_rom.i_col\[4\] vssd1 vssd1
+ vccd1 vccd1 _03973_ sky130_fd_sc_hd__and3_1
XFILLER_122_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17800_ _09668_ _09552_ _09973_ _08802_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__o22a_1
XFILLER_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18780_ rbzero.wall_tracer.trackDistY\[-2\] rbzero.wall_tracer.stepDistY\[-2\] vssd1
+ vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__nor2_1
X_15992_ _08634_ _08636_ vssd1 vssd1 vccd1 vccd1 _08637_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17731_ _10294_ _10184_ _10185_ vssd1 vssd1 vccd1 vccd1 _10296_ sky130_fd_sc_hd__or3_1
XFILLER_134_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14943_ rbzero.wall_tracer.trackDistY\[6\] rbzero.wall_tracer.trackDistX\[6\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__mux2_1
XFILLER_169_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17662_ _10070_ _10079_ _10226_ vssd1 vssd1 vccd1 vccd1 _10227_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14874_ _07452_ _07451_ _05892_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__mux2_1
XFILLER_29_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19401_ _02873_ _02884_ _02885_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__or3_1
X_16613_ _09254_ _09255_ vssd1 vssd1 vccd1 vccd1 _09256_ sky130_fd_sc_hd__xnor2_1
X_13825_ _06561_ _06276_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__xor2_2
X_17593_ _10156_ _10158_ vssd1 vssd1 vccd1 vccd1 _10159_ sky130_fd_sc_hd__xor2_1
XFILLER_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16544_ _09186_ _09187_ vssd1 vssd1 vccd1 vccd1 _09188_ sky130_fd_sc_hd__xnor2_4
X_19332_ rbzero.pov.spi_done rbzero.pov.ready _02730_ _02823_ vssd1 vssd1 vccd1 vccd1
+ _00804_ sky130_fd_sc_hd__o211a_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13756_ _06491_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__nor2_1
XFILLER_90_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10968_ rbzero.tex_b1\[8\] rbzero.tex_b1\[9\] _03828_ vssd1 vssd1 vccd1 vccd1 _03832_
+ sky130_fd_sc_hd__mux2_1
X_12707_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[9\] _05446_
+ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__a21bo_1
X_16475_ _08284_ _08177_ vssd1 vssd1 vccd1 vccd1 _09119_ sky130_fd_sc_hd__nor2_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19263_ _02785_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13687_ _06422_ _06423_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__and2_1
X_10899_ rbzero.tex_b1\[41\] rbzero.tex_b1\[42\] _03795_ vssd1 vssd1 vccd1 vccd1 _03796_
+ sky130_fd_sc_hd__mux2_1
XFILLER_176_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18214_ _01908_ _01914_ rbzero.wall_tracer.trackDistX\[6\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00595_ sky130_fd_sc_hd__o2bb2a_1
X_15426_ _08070_ rbzero.debug_overlay.playerY\[-3\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _08071_ sky130_fd_sc_hd__mux2_1
XFILLER_54_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19194_ rbzero.spi_registers.new_sky\[1\] rbzero.color_sky\[1\] _02740_ vssd1 vssd1
+ vccd1 vccd1 _02743_ sky130_fd_sc_hd__mux2_1
X_12638_ _05389_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__inv_2
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18145_ _01844_ _01845_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__nand2_1
XFILLER_157_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15357_ _07904_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__clkbuf_4
X_12569_ _05321_ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__and2_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14308_ _06134_ _06662_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__nor2_1
XFILLER_89_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18076_ _01653_ _01654_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__nor2_1
X_15288_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__buf_4
XFILLER_144_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17027_ _09665_ _09666_ vssd1 vssd1 vccd1 vccd1 _09667_ sky130_fd_sc_hd__nand2_1
XFILLER_160_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14239_ _06970_ _06975_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__xor2_1
XFILLER_98_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18978_ _02619_ vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__clkbuf_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _01613_ _01631_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__xor2_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20940_ clknet_leaf_9_i_clk _00709_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_93_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19640__90 clknet_1_0__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__inv_2
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20871_ clknet_leaf_94_i_clk _00640_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20243__263 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__inv_2
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21423_ net344 _01192_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21354_ net275 _01123_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20305_ clknet_1_1__leaf__03309_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__buf_1
XFILLER_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21285_ clknet_leaf_38_i_clk _01054_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_151_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20326__338 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__inv_2
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _04230_ _04711_ _04715_ _04242_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__a211o_1
XFILLER_45_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _04646_ _04647_ _04217_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__mux2_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _06345_ _06346_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__nor2_1
XFILLER_38_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10822_ _03755_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__clkbuf_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _07203_ _07210_ _07154_ vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__a21oi_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13541_ _06193_ _06231_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__xor2_1
X_10753_ _03719_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16260_ _08902_ _08904_ vssd1 vssd1 vccd1 vccd1 _08905_ sky130_fd_sc_hd__nor2_1
XFILLER_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13472_ _06168_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__xnor2_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10684_ rbzero.tex_g1\[15\] rbzero.tex_g1\[16\] _03680_ vssd1 vssd1 vccd1 vccd1 _03683_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15211_ _04034_ _07861_ _07862_ _07718_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__o31a_1
X_12423_ _05187_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__buf_2
XFILLER_200_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16191_ _08815_ _08835_ vssd1 vssd1 vccd1 vccd1 _08836_ sky130_fd_sc_hd__xor2_1
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15142_ _07786_ _07789_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__and2_1
X_12354_ _05101_ _05120_ _05121_ net31 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__o211a_1
XFILLER_127_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20071__108 clknet_1_0__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__inv_2
X_11305_ rbzero.traced_texVinit\[1\] rbzero.texV\[1\] rbzero.texV\[0\] rbzero.traced_texVinit\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__o211a_1
X_15073_ _07732_ _07733_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__xnor2_1
X_19950_ _03241_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__buf_2
X_12285_ net46 _05046_ _05049_ _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__a22o_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18901_ rbzero.spi_registers.spi_counter\[3\] _02564_ _02570_ vssd1 vssd1 vccd1 vccd1
+ _02571_ sky130_fd_sc_hd__o21a_1
X_14024_ _05752_ _06658_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__nand2_2
X_11236_ gpout0.hpos\[9\] _04009_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__and2_2
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19881_ _03188_ _03186_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__nor2_1
XFILLER_150_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18832_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.stepDistY\[5\] vssd1
+ vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__or2_1
X_11167_ rbzero.otherx\[1\] rbzero.map_rom.f3 vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__xor2_1
XFILLER_68_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18763_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.stepDistY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__nor2_1
XFILLER_110_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15975_ _08609_ _08611_ vssd1 vssd1 vccd1 vccd1 _08620_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19614__68 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__inv_2
X_11098_ rbzero.tex_b0\[11\] rbzero.tex_b0\[10\] _03898_ vssd1 vssd1 vccd1 vccd1 _03900_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17714_ _10109_ _10151_ _10278_ vssd1 vssd1 vccd1 vccd1 _10279_ sky130_fd_sc_hd__a21bo_1
XFILLER_36_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14926_ rbzero.wall_tracer.visualWallDist\[0\] _07618_ vssd1 vssd1 vccd1 vccd1 _07627_
+ sky130_fd_sc_hd__or2_1
X_18694_ _09889_ _02388_ _02389_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__or3b_1
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17645_ _09096_ _09359_ _10060_ _10059_ vssd1 vssd1 vccd1 vccd1 _10210_ sky130_fd_sc_hd__o31a_1
XFILLER_24_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14857_ _07468_ _07574_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__nand2b_4
XFILLER_17_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _06490_ _06493_ _06494_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__or3_1
XFILLER_51_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17576_ _10137_ _10140_ _10141_ vssd1 vssd1 vccd1 vccd1 _10142_ sky130_fd_sc_hd__and3_1
X_14788_ _05884_ _07477_ _07419_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__or3_1
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19315_ rbzero.spi_registers.new_vshift\[0\] rbzero.spi_registers.spi_buffer\[0\]
+ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__mux2_1
X_16527_ _09169_ _09170_ vssd1 vssd1 vccd1 vccd1 _09171_ sky130_fd_sc_hd__nand2_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13739_ _06045_ _06009_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__nor2_1
XFILLER_56_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19246_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_sky\[1\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__mux2_1
XFILLER_91_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16458_ _09100_ _09101_ vssd1 vssd1 vccd1 vccd1 _09102_ sky130_fd_sc_hd__xnor2_1
XFILLER_143_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15409_ _08053_ vssd1 vssd1 vccd1 vccd1 _08054_ sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__04835_ clknet_0__04835_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__04835_
+ sky130_fd_sc_hd__clkbuf_16
X_16389_ _09032_ _09033_ vssd1 vssd1 vccd1 vccd1 _09034_ sky130_fd_sc_hd__nand2_1
X_19177_ rbzero.spi_registers.got_new_leak _02711_ vssd1 vssd1 vccd1 vccd1 _02733_
+ sky130_fd_sc_hd__nand2_1
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18128_ _01827_ _01828_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__xnor2_1
XFILLER_157_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20273__289 clknet_1_1__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__inv_2
X_18059_ _01757_ _01758_ _01759_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a21o_1
XFILLER_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21070_ net160 _00839_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20021_ _04990_ _04989_ _03258_ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__or4_1
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20167__194 clknet_1_0__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__inv_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20923_ clknet_leaf_22_i_clk _00692_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20384__10 clknet_1_0__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__inv_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20854_ clknet_leaf_51_i_clk _00623_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20785_ clknet_leaf_27_i_clk _00554_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_57_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21406_ net327 _01175_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[49\] sky130_fd_sc_hd__dfxtp_1
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21337_ net258 _01106_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12070_ _04840_ _04666_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__nand2_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21268_ clknet_leaf_89_i_clk _01037_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneY\[-9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11021_ _03859_ vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__clkbuf_1
X_21199_ clknet_leaf_99_i_clk _00968_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi sky130_fd_sc_hd__dfxtp_1
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _08337_ _08347_ vssd1 vssd1 vccd1 vccd1 _08405_ sky130_fd_sc_hd__xnor2_1
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12972_ _05563_ _05566_ _05600_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__and3_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _07375_ _07447_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__or2_1
X_11923_ _04241_ _04690_ _04698_ _04207_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__o211a_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _08059_ _08335_ vssd1 vssd1 vccd1 vccd1 _08336_ sky130_fd_sc_hd__nor2_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _07601_ _09995_ _09996_ vssd1 vssd1 vccd1 vccd1 _09997_ sky130_fd_sc_hd__mux2_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14642_ _07378_ _07349_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__nand2_1
XFILLER_79_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ rbzero.tex_g1\[13\] rbzero.tex_g1\[12\] _04337_ vssd1 vssd1 vccd1 vccd1 _04631_
+ sky130_fd_sc_hd__mux2_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _03746_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__clkbuf_1
X_17361_ _09243_ _09029_ _09164_ _09096_ vssd1 vssd1 vccd1 vccd1 _09928_ sky130_fd_sc_hd__o22ai_1
X_14573_ _07305_ _07093_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__xnor2_1
XFILLER_198_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11785_ _04560_ _04561_ _04562_ _04304_ _04253_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__o221a_1
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19100_ _02683_ vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13524_ _06259_ _06260_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__nor2_1
X_16312_ _08550_ _08616_ _08673_ _08955_ _08956_ vssd1 vssd1 vccd1 vccd1 _08957_ sky130_fd_sc_hd__o221ai_4
XFILLER_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10736_ rbzero.tex_g0\[55\] rbzero.tex_g0\[54\] _03706_ vssd1 vssd1 vccd1 vccd1 _03710_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17292_ rbzero.wall_tracer.trackDistX\[-5\] rbzero.wall_tracer.stepDistX\[-5\] vssd1
+ vssd1 vccd1 vccd1 _09864_ sky130_fd_sc_hd__or2_1
XFILLER_203_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16243_ _08871_ _08887_ vssd1 vssd1 vccd1 vccd1 _08888_ sky130_fd_sc_hd__nand2_1
X_19031_ rbzero.pov.spi_buffer\[47\] rbzero.pov.ready_buffer\[47\] _02638_ vssd1 vssd1
+ vccd1 vccd1 _02647_ sky130_fd_sc_hd__mux2_1
X_13455_ _06189_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__xnor2_1
XFILLER_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ rbzero.tex_g1\[23\] rbzero.tex_g1\[24\] _03669_ vssd1 vssd1 vccd1 vccd1 _03674_
+ sky130_fd_sc_hd__mux2_1
XFILLER_173_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12406_ _04883_ _04884_ _04886_ _04887_ _05143_ net34 vssd1 vssd1 vccd1 vccd1 _05173_
+ sky130_fd_sc_hd__mux4_1
XFILLER_127_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16174_ _08816_ _08075_ _08817_ _08784_ vssd1 vssd1 vccd1 vccd1 _08819_ sky130_fd_sc_hd__o22a_1
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13386_ _06041_ _05991_ _05940_ _06078_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__o22ai_1
XFILLER_182_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10598_ _03637_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15125_ _07782_ vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__clkbuf_1
X_12337_ net46 _05103_ _05104_ _05099_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15056_ rbzero.wall_tracer.rayAddendX\[-3\] _07717_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07719_ sky130_fd_sc_hd__mux2_1
X_19933_ rbzero.debug_overlay.playerY\[3\] _03223_ _02822_ vssd1 vssd1 vccd1 vccd1
+ _03228_ sky130_fd_sc_hd__a21o_1
XFILLER_114_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12268_ _04886_ _04887_ _05021_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__mux2_1
XFILLER_142_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14007_ _06666_ _06708_ _06742_ _06743_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__o31ai_2
X_11219_ gpout0.hpos\[6\] vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__clkbuf_4
X_19864_ rbzero.debug_overlay.playerX\[1\] _03143_ _03174_ _03175_ vssd1 vssd1 vccd1
+ vccd1 _00984_ sky130_fd_sc_hd__a211o_1
X_12199_ net17 net18 vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__nand2_1
X_18815_ _05532_ _02494_ _02495_ _02399_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__o31a_1
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20309__322 clknet_1_0__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__inv_2
X_19795_ _03126_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18746_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.stepDistY\[-6\] vssd1
+ vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__03295_ clknet_0__03295_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03295_
+ sky130_fd_sc_hd__clkbuf_16
X_15958_ _08588_ _08600_ vssd1 vssd1 vccd1 vccd1 _08603_ sky130_fd_sc_hd__nor2_1
XFILLER_49_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14909_ rbzero.wall_tracer.trackDistY\[-4\] rbzero.wall_tracer.trackDistX\[-4\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__mux2_1
XFILLER_184_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18677_ _02368_ _02372_ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15889_ _08531_ _08532_ _08533_ vssd1 vssd1 vccd1 vccd1 _08534_ sky130_fd_sc_hd__a21oi_1
XFILLER_24_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17628_ _10085_ _10187_ _10191_ vssd1 vssd1 vccd1 vccd1 _10193_ sky130_fd_sc_hd__and3_1
XFILLER_197_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17559_ _08747_ _09700_ vssd1 vssd1 vccd1 vccd1 _10125_ sky130_fd_sc_hd__nor2_1
XFILLER_176_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20570_ gpout0.clk_div\[0\] gpout0.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__nand2_1
XFILLER_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19229_ rbzero.spi_registers.new_vshift\[1\] _02763_ vssd1 vssd1 vccd1 vccd1 _02766_
+ sky130_fd_sc_hd__or2_1
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20355__364 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__inv_2
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21122_ net212 _00891_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21053_ clknet_leaf_99_i_clk _00822_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20004_ rbzero.pov.ready_buffer\[8\] _03239_ _03242_ rbzero.debug_overlay.vplaneY\[-1\]
+ _02730_ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__o221a_1
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20906_ clknet_leaf_91_i_clk _00675_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20837_ clknet_leaf_53_i_clk _00606_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11570_ rbzero.tex_r1\[3\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__and3_1
XFILLER_126_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20768_ clknet_leaf_45_i_clk _00537_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10521_ rbzero.tex_r0\[29\] rbzero.tex_r0\[28\] _03591_ vssd1 vssd1 vccd1 vccd1 _03597_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20699_ clknet_leaf_49_i_clk _00483_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_149_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _05962_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__nand2_1
XFILLER_7_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10452_ rbzero.tex_r0\[62\] rbzero.tex_r0\[61\] _03558_ vssd1 vssd1 vccd1 vccd1 _03561_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13171_ _05884_ _05859_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__or2_1
X_10383_ _03522_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_151_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12122_ _04885_ _04888_ _04889_ _04893_ net4 net3 vssd1 vssd1 vccd1 vccd1 _04894_
+ sky130_fd_sc_hd__mux4_2
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16930_ _09559_ _09570_ vssd1 vssd1 vccd1 vccd1 _09571_ sky130_fd_sc_hd__xnor2_2
X_12053_ rbzero.row_render.side _04821_ _04826_ _04814_ _04820_ vssd1 vssd1 vccd1
+ vccd1 _04827_ sky130_fd_sc_hd__o221ai_1
XFILLER_46_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11004_ _03850_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_46_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16861_ _09243_ _08159_ _08150_ _09245_ vssd1 vssd1 vccd1 vccd1 _09502_ sky130_fd_sc_hd__o22a_1
XFILLER_133_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18600_ _02179_ _02182_ _02295_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__and3_1
X_15812_ _08025_ _08013_ vssd1 vssd1 vccd1 vccd1 _08457_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16792_ _09429_ _09433_ _05209_ vssd1 vssd1 vccd1 vccd1 _09434_ sky130_fd_sc_hd__a21o_2
XFILLER_206_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18531_ rbzero.wall_tracer.trackDistX\[9\] rbzero.wall_tracer.stepDistX\[9\] vssd1
+ vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__or2_1
X_15743_ _08386_ _08387_ vssd1 vssd1 vccd1 vccd1 _08388_ sky130_fd_sc_hd__xnor2_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _05642_ _05645_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__or2_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _04332_ _04677_ _04681_ _04142_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a211o_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18462_ _02143_ _02159_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__xnor2_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15674_ _08263_ _08264_ _08307_ vssd1 vssd1 vccd1 vccd1 _08319_ sky130_fd_sc_hd__and3_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _05609_ _05619_ _05622_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__or3_1
XFILLER_93_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _08284_ _09540_ vssd1 vssd1 vccd1 vccd1 _09980_ sky130_fd_sc_hd__nor2_2
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11837_ rbzero.tex_g1\[45\] rbzero.tex_g1\[44\] _04337_ vssd1 vssd1 vccd1 vccd1 _04614_
+ sky130_fd_sc_hd__mux2_1
X_14625_ _07357_ _07361_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__or2_1
X_18393_ _02086_ _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__xnor2_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17344_ _08335_ _09359_ _09910_ _09624_ vssd1 vssd1 vccd1 vccd1 _09911_ sky130_fd_sc_hd__o31a_1
X_14556_ _07286_ _07292_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__nor2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _04542_ _04545_ _04208_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__mux2_1
XFILLER_186_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10719_ rbzero.tex_g0\[63\] rbzero.tex_g0\[62\] _03624_ vssd1 vssd1 vccd1 vccd1 _03701_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13507_ _05983_ _05940_ _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__or3_1
XFILLER_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14487_ _07177_ _07009_ _07223_ _07065_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__a22o_1
X_17275_ _09846_ _09847_ _09848_ vssd1 vssd1 vccd1 vccd1 _09849_ sky130_fd_sc_hd__and3_1
X_11699_ rbzero.debug_overlay.vplaneY\[10\] _04453_ _04474_ _04477_ vssd1 vssd1 vccd1
+ vccd1 _04478_ sky130_fd_sc_hd__a211o_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19014_ _02594_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__buf_4
X_16226_ _08870_ vssd1 vssd1 vccd1 vccd1 _08871_ sky130_fd_sc_hd__inv_2
X_13438_ _05998_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__or2_1
X_16157_ _08111_ vssd1 vssd1 vccd1 vccd1 _08802_ sky130_fd_sc_hd__buf_4
X_13369_ _06099_ _06102_ _06105_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__nand3_1
XFILLER_182_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15108_ _07749_ _07766_ vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__xnor2_1
X_16088_ _08284_ _08128_ _08727_ _08732_ vssd1 vssd1 vccd1 vccd1 _08733_ sky130_fd_sc_hd__o31ai_2
XFILLER_170_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15039_ _03913_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__clkbuf_4
XFILLER_69_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19916_ _08089_ _03164_ _03193_ _03214_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__a211oi_1
XFILLER_69_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19847_ rbzero.pov.ready_buffer\[66\] _08077_ _03146_ vssd1 vssd1 vccd1 vccd1 _03162_
+ sky130_fd_sc_hd__mux2_1
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19778_ rbzero.pov.spi_buffer\[62\] rbzero.pov.spi_buffer\[63\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03118_ sky130_fd_sc_hd__mux2_1
XFILLER_95_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18729_ _02420_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20622_ clknet_leaf_15_i_clk _00406_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.mapY\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_189_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20279__295 clknet_1_0__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__inv_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20553_ _03436_ _03439_ _03440_ _09748_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__a31o_1
XFILLER_193_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20484_ rbzero.traced_texa\[0\] rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 _03384_
+ sky130_fd_sc_hd__nand2_1
XFILLER_138_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21105_ net195 _00874_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21036_ clknet_leaf_77_i_clk _00805_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12740_ _05486_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__xnor2_2
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ rbzero.debug_overlay.facingX\[-4\] rbzero.wall_tracer.rayAddendX\[4\] vssd1
+ vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__nor2_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14410_ _07120_ _07126_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__or2_1
XFILLER_70_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11622_ rbzero.tex_r1\[33\] rbzero.tex_r1\[32\] _04392_ vssd1 vssd1 vccd1 vccd1 _04401_
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15390_ _08034_ vssd1 vssd1 vccd1 vccd1 _08035_ sky130_fd_sc_hd__clkbuf_4
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14341_ _07017_ _07019_ _06774_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__o21ai_1
XFILLER_204_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ _04208_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__buf_4
XFILLER_195_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10504_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _03580_ vssd1 vssd1 vccd1 vccd1 _03588_
+ sky130_fd_sc_hd__mux2_1
X_17060_ _08816_ _09699_ vssd1 vssd1 vccd1 vccd1 _09700_ sky130_fd_sc_hd__or2_2
X_14272_ _06675_ _06740_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__nor2_1
XFILLER_184_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11484_ rbzero.tex_r0\[37\] rbzero.tex_r0\[36\] _04263_ vssd1 vssd1 vccd1 vccd1 _04264_
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16011_ _08634_ _08636_ _08655_ vssd1 vssd1 vccd1 vccd1 _08656_ sky130_fd_sc_hd__a21bo_1
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03298_ clknet_0__03298_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03298_
+ sky130_fd_sc_hd__clkbuf_16
X_13223_ _05901_ _05831_ _05956_ _05959_ _05871_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a2111o_1
X_10435_ rbzero.tex_r1\[3\] rbzero.tex_r1\[4\] _03549_ vssd1 vssd1 vccd1 vccd1 _03550_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13154_ _05872_ _05890_ _05826_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__mux2_1
X_10366_ _03513_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12105_ net5 _04850_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__or2_1
XFILLER_135_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17962_ _01546_ _01442_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__or2b_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13085_ _05814_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__or2_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19701_ _03077_ vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__clkbuf_1
X_12036_ _04317_ _04163_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__nor2_1
X_16913_ rbzero.wall_tracer.stepDistX\[7\] vssd1 vssd1 vccd1 vccd1 _09554_ sky130_fd_sc_hd__inv_2
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17893_ _01594_ _01595_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__03301_ _03301_ vssd1 vssd1 vccd1 vccd1 clknet_0__03301_ sky130_fd_sc_hd__clkbuf_16
X_16844_ _08160_ _09480_ _09484_ _08162_ vssd1 vssd1 vccd1 vccd1 _09485_ sky130_fd_sc_hd__o22ai_1
XFILLER_66_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19563_ _03031_ _03020_ _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__and3b_1
X_16775_ _09416_ vssd1 vssd1 vccd1 vccd1 _09417_ sky130_fd_sc_hd__clkbuf_4
XFILLER_168_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13987_ _06067_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__clkbuf_4
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18514_ _02205_ _02206_ _02210_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__and3_1
XFILLER_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15726_ _08327_ _08370_ vssd1 vssd1 vccd1 vccd1 _08371_ sky130_fd_sc_hd__xnor2_2
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19494_ _02904_ rbzero.wall_tracer.rayAddendY\[7\] vssd1 vssd1 vccd1 vccd1 _02973_
+ sky130_fd_sc_hd__nand2_1
X_12938_ _05659_ _05603_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__nand2_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18445_ _02044_ _02052_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__a21o_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ _08300_ _08301_ vssd1 vssd1 vccd1 vccd1 _08302_ sky130_fd_sc_hd__xnor2_1
X_12869_ _05603_ _05605_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__nand2_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ _07330_ _07342_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__xnor2_1
X_18376_ _02073_ _02074_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__xor2_1
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15588_ _08218_ _08208_ _08232_ vssd1 vssd1 vccd1 vccd1 _08233_ sky130_fd_sc_hd__a21oi_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17327_ rbzero.wall_tracer.trackDistX\[-2\] _09817_ _09888_ _09895_ vssd1 vssd1 vccd1
+ vccd1 _00587_ sky130_fd_sc_hd__o22a_1
XFILLER_119_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14539_ _07274_ _07275_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__nor2_1
XFILLER_174_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17258_ _09830_ _09831_ _09832_ vssd1 vssd1 vccd1 vccd1 _09834_ sky130_fd_sc_hd__a21oi_1
XFILLER_179_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16209_ _08519_ _08053_ vssd1 vssd1 vccd1 vccd1 _08854_ sky130_fd_sc_hd__nor2_1
X_17189_ rbzero.wall_tracer.mapX\[6\] _05512_ vssd1 vssd1 vccd1 vccd1 _09774_ sky130_fd_sc_hd__xor2_1
XFILLER_108_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21654_ clknet_leaf_37_i_clk _01423_ vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20605_ gpout3.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__nor2_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21585_ net506 _01354_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xtop_ew_algofoogle_77 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_77/HI o_rgb[5] sky130_fd_sc_hd__conb_1
X_20536_ rbzero.traced_texa\[7\] rbzero.texV\[7\] _03427_ vssd1 vssd1 vccd1 vccd1
+ _03428_ sky130_fd_sc_hd__o21ai_1
Xtop_ew_algofoogle_88 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_88/HI o_rgb[20] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_99 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_99/HI zeros[9] sky130_fd_sc_hd__conb_1
XFILLER_181_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20467_ _03367_ _03368_ _03369_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__a21o_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13910_ _05752_ _05989_ _06053_ _06624_ _06646_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__a41o_1
X_21019_ clknet_leaf_9_i_clk _00788_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14890_ rbzero.wall_tracer.visualWallDist\[-10\] vssd1 vssd1 vccd1 vccd1 _07601_
+ sky130_fd_sc_hd__buf_4
XFILLER_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13841_ _06576_ _06577_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__and2_1
XFILLER_75_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16560_ _05194_ _09202_ _09203_ _07642_ vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__o211a_1
X_13772_ _06508_ _06481_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__xnor2_1
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10984_ rbzero.tex_b1\[0\] rbzero.tex_b1\[1\] _03482_ vssd1 vssd1 vccd1 vccd1 _03840_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15511_ _08056_ _08063_ vssd1 vssd1 vccd1 vccd1 _08156_ sky130_fd_sc_hd__and2_1
X_12723_ _05422_ _05429_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__and2b_1
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16491_ _09133_ _09134_ vssd1 vssd1 vccd1 vccd1 _09135_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18230_ _01874_ _01858_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__or2b_1
X_15442_ _08076_ _08085_ vssd1 vssd1 vccd1 vccd1 _08087_ sky130_fd_sc_hd__nand2_1
X_12654_ _05397_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__clkbuf_4
XFILLER_203_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ rbzero.tex_r1\[49\] rbzero.tex_r1\[48\] _04338_ vssd1 vssd1 vccd1 vccd1 _04384_
+ sky130_fd_sc_hd__mux2_1
X_18161_ _01859_ _01861_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__nand2_1
X_12585_ _05296_ _05297_ _05337_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__nand3b_1
X_15373_ _07903_ rbzero.wall_tracer.stepDistY\[-7\] _05195_ vssd1 vssd1 vccd1 vccd1
+ _08018_ sky130_fd_sc_hd__a21o_1
XFILLER_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17112_ _09749_ vssd1 vssd1 vccd1 vccd1 _09750_ sky130_fd_sc_hd__clkbuf_4
XFILLER_128_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11536_ gpout0.vpos\[5\] gpout0.vpos\[3\] vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__nand2_1
X_14324_ _07060_ _06843_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__nand2_1
XFILLER_184_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18092_ rbzero.wall_tracer.trackDistX\[5\] rbzero.wall_tracer.stepDistX\[5\] vssd1
+ vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__nand2_1
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17043_ _09553_ _09557_ _09556_ vssd1 vssd1 vccd1 vccd1 _09683_ sky130_fd_sc_hd__a21bo_1
X_14255_ _06962_ _06984_ _06988_ _06951_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__o22a_1
XFILLER_7_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11467_ _04139_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__buf_4
XFILLER_125_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _05846_ _05940_ _05942_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__or3_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10418_ rbzero.tex_r1\[11\] rbzero.tex_r1\[12\] _03538_ vssd1 vssd1 vccd1 vccd1 _03541_
+ sky130_fd_sc_hd__mux2_1
X_14186_ _06921_ _06922_ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__xnor2_1
X_11398_ rbzero.row_render.size\[8\] rbzero.row_render.size\[7\] _04152_ vssd1 vssd1
+ vccd1 vccd1 _04178_ sky130_fd_sc_hd__nor3_1
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _05778_ _05872_ _05873_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__o21a_1
X_10349_ _03504_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__clkbuf_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18994_ rbzero.pov.spi_buffer\[29\] rbzero.pov.ready_buffer\[29\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02628_ sky130_fd_sc_hd__mux2_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _01643_ _01644_ _01646_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a21o_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _05721_ _05734_ _05796_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__mux2_1
XFILLER_79_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12019_ _04379_ _04791_ _04792_ _04793_ _04209_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__o221a_1
X_17876_ _09096_ _09703_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__nand2_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19615_ clknet_1_1__leaf__03037_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__buf_1
X_16827_ _09082_ _09467_ _05194_ vssd1 vssd1 vccd1 vccd1 _09469_ sky130_fd_sc_hd__a21o_1
XFILLER_54_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19546_ rbzero.pov.ss_buffer\[1\] _03555_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__nor2_2
XFILLER_65_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16758_ _09252_ _09394_ _09399_ vssd1 vssd1 vccd1 vccd1 _09400_ sky130_fd_sc_hd__a21oi_1
XFILLER_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15709_ _08352_ _08353_ vssd1 vssd1 vccd1 vccd1 _08354_ sky130_fd_sc_hd__nand2_1
X_19477_ _02941_ _02944_ _02957_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__o21a_1
X_16689_ rbzero.debug_overlay.playerY\[-4\] vssd1 vssd1 vccd1 vccd1 _09332_ sky130_fd_sc_hd__inv_2
XFILLER_34_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18428_ _02125_ _02126_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__nand2_1
XFILLER_179_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18359_ _02056_ _02057_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__nor2_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21370_ net291 _01139_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20183_ clknet_1_0__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__buf_1
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20220__242 clknet_1_1__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__inv_2
XFILLER_185_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21637_ clknet_leaf_41_i_clk _01406_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12370_ _04738_ _05086_ _05098_ _05137_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__o2bb2a_2
XFILLER_201_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21568_ net489 _01337_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11321_ _04060_ _04063_ _04100_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__o21ba_1
XFILLER_10_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20519_ _03406_ _03407_ _03408_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__o21ai_1
XFILLER_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21499_ net420 _01268_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[14\] sky130_fd_sc_hd__dfxtp_1
X_14040_ _06776_ _06658_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__nor2_1
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11252_ _04033_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__buf_4
XFILLER_84_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11183_ rbzero.map_rom.d6 _03942_ _03933_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_
+ sky130_fd_sc_hd__and4_1
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15991_ _08635_ _08561_ vssd1 vssd1 vccd1 vccd1 _08636_ sky130_fd_sc_hd__xnor2_1
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17730_ _10184_ _10185_ _10294_ vssd1 vssd1 vccd1 vccd1 _10295_ sky130_fd_sc_hd__o21a_1
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14942_ _07621_ _07636_ _07637_ _07620_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__o211a_1
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17661_ _10071_ _09961_ _10078_ vssd1 vssd1 vccd1 vccd1 _10226_ sky130_fd_sc_hd__a21oi_1
X_14873_ _07587_ vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19400_ _02884_ _02885_ _02873_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__o21ai_1
X_16612_ _07996_ _09103_ vssd1 vssd1 vccd1 vccd1 _09255_ sky130_fd_sc_hd__or2_1
X_13824_ _06193_ _06231_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__nand2_1
XFILLER_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17592_ _09955_ _10014_ _10157_ vssd1 vssd1 vccd1 vccd1 _10158_ sky130_fd_sc_hd__a21boi_1
XFILLER_16_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20303__317 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__inv_2
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19331_ _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__clkbuf_4
X_16543_ _09046_ _09048_ _09045_ vssd1 vssd1 vccd1 vccd1 _09187_ sky130_fd_sc_hd__a21boi_4
X_13755_ _06467_ _06489_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__xor2_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10967_ _03831_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ _05450_ _05453_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__xnor2_2
X_19262_ rbzero.spi_registers.spi_buffer\[1\] rbzero.spi_registers.new_floor\[1\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__mux2_1
XFILLER_149_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16474_ _08178_ _09117_ _08972_ _08973_ vssd1 vssd1 vccd1 vccd1 _09118_ sky130_fd_sc_hd__o31ai_2
XFILLER_31_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13686_ _06336_ _06375_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__xor2_1
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10898_ _03646_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__clkbuf_4
XFILLER_188_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18213_ _01912_ _01913_ _09780_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__a21oi_1
XFILLER_54_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15425_ _08029_ _08069_ vssd1 vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__and2_1
XFILLER_19_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19193_ rbzero.color_sky\[0\] _02740_ _02742_ vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__a21o_1
X_12637_ rbzero.map_rom.a6 _05374_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__and2_1
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18144_ _10239_ _08423_ _01843_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__o21ai_1
XFILLER_156_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12568_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] vssd1
+ vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__nand2_1
X_15356_ _07999_ _08000_ _05496_ vssd1 vssd1 vccd1 vccd1 _08001_ sky130_fd_sc_hd__mux2_2
XFILLER_200_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11519_ rbzero.tex_r0\[27\] rbzero.tex_r0\[26\] _04263_ vssd1 vssd1 vccd1 vccd1 _04299_
+ sky130_fd_sc_hd__mux2_1
XFILLER_157_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14307_ _07005_ _06731_ _06700_ _07004_ _07003_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__o32ai_4
XFILLER_89_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18075_ _01775_ _01776_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__or2_1
XFILLER_141_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15287_ _07931_ vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__clkbuf_4
XFILLER_89_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12499_ rbzero.wall_tracer.trackDistY\[2\] vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__inv_2
XFILLER_156_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17026_ _09661_ _08047_ _09662_ _09664_ vssd1 vssd1 vccd1 vccd1 _09666_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_172_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14238_ _06935_ _06963_ _06972_ _06974_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__a31o_1
XFILLER_153_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14169_ _06904_ _06903_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__and2b_1
XFILLER_124_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ rbzero.pov.spi_buffer\[21\] rbzero.pov.ready_buffer\[21\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02619_ sky130_fd_sc_hd__mux2_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _01615_ _01630_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__xor2_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17859_ _01491_ _01455_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__or2b_1
XFILLER_27_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20870_ clknet_leaf_93_i_clk _00639_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19529_ _02994_ _02995_ _02998_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__mux2_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_1_i_clk clknet_1_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1_1_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_194_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21422_ net343 _01191_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21353_ net274 _01122_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21284_ clknet_leaf_38_i_clk _01053_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ rbzero.tex_g1\[17\] rbzero.tex_g1\[16\] _04211_ vssd1 vssd1 vccd1 vccd1 _04647_
+ sky130_fd_sc_hd__mux2_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ rbzero.tex_g0\[15\] rbzero.tex_g0\[14\] _03751_ vssd1 vssd1 vccd1 vccd1 _03755_
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20999_ clknet_leaf_13_i_clk _00768_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10752_ rbzero.tex_g0\[48\] rbzero.tex_g0\[47\] _03718_ vssd1 vssd1 vccd1 vccd1 _03719_
+ sky130_fd_sc_hd__mux2_1
X_13540_ _06193_ _06231_ _06276_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__and3_1
XFILLER_38_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13471_ _06199_ _06207_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__xnor2_1
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ _03682_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15210_ _07850_ _07854_ _07860_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__a21oi_1
X_12422_ net71 rbzero.wall_tracer.state\[9\] _03480_ vssd1 vssd1 vccd1 vccd1 _05187_
+ sky130_fd_sc_hd__and3_1
X_16190_ _08827_ _08833_ _08834_ vssd1 vssd1 vccd1 vccd1 _08835_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12353_ net29 _05094_ net30 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__o21ai_1
X_15141_ _07785_ rbzero.wall_tracer.rayAddendX\[4\] vssd1 vssd1 vccd1 vccd1 _07797_
+ sky130_fd_sc_hd__xor2_1
XFILLER_5_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11304_ rbzero.texV\[3\] _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__xor2_1
X_15072_ _07721_ _07724_ _07722_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__a21bo_1
X_12284_ _04867_ _05034_ _05027_ net47 vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__a31o_1
XFILLER_126_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18900_ rbzero.spi_registers.spi_counter\[1\] _02569_ vssd1 vssd1 vccd1 vccd1 _02570_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14023_ _06758_ _06759_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__nand2_4
XFILLER_135_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11235_ _04015_ _04019_ _03914_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__a21oi_1
X_19880_ rbzero.debug_overlay.playerX\[5\] vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__inv_2
XFILLER_175_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18831_ _02509_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__clkbuf_1
X_11166_ _03915_ _03918_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__o21a_1
XFILLER_84_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18762_ _02449_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11097_ _03899_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__clkbuf_1
X_15974_ _08584_ _08618_ vssd1 vssd1 vccd1 vccd1 _08619_ sky130_fd_sc_hd__xnor2_4
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17713_ _10147_ _10150_ vssd1 vssd1 vccd1 vccd1 _10278_ sky130_fd_sc_hd__or2b_1
X_14925_ rbzero.wall_tracer.trackDistY\[0\] rbzero.wall_tracer.trackDistX\[0\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__mux2_1
X_18693_ _02310_ _02313_ _02387_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__or3_1
XFILLER_64_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ _10207_ _10208_ vssd1 vssd1 vccd1 vccd1 _10209_ sky130_fd_sc_hd__xnor2_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14856_ _07433_ _07374_ _07573_ _07394_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__o211ai_4
XFILLER_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13807_ _06505_ _06524_ _06525_ _06543_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__o211a_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17575_ _08872_ _10139_ _08266_ _09989_ vssd1 vssd1 vccd1 vccd1 _10141_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14787_ _05884_ _07516_ _07518_ _05800_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__a211o_1
XFILLER_95_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11999_ _04772_ _04773_ _04225_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__mux2_1
XFILLER_182_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19314_ _02812_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__clkbuf_4
X_16526_ _08112_ _08150_ _08331_ _08417_ vssd1 vssd1 vccd1 vccd1 _09170_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13738_ _05846_ _05823_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__nor2_1
XFILLER_108_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19245_ _02775_ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__clkbuf_1
XFILLER_182_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16457_ _07932_ _08097_ vssd1 vssd1 vccd1 vccd1 _09101_ sky130_fd_sc_hd__or2_1
X_13669_ _05856_ _05877_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__nand2_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15408_ _07903_ _08048_ _08051_ _08052_ _05196_ vssd1 vssd1 vccd1 vccd1 _08053_ sky130_fd_sc_hd__o311a_4
X_19176_ _02731_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__clkbuf_2
X_16388_ _08053_ _08158_ _08418_ _08039_ vssd1 vssd1 vccd1 vccd1 _09033_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18127_ _10094_ _09027_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__nor2_1
X_15339_ rbzero.wall_tracer.visualWallDist\[-8\] _07983_ _07903_ vssd1 vssd1 vccd1
+ vccd1 _07984_ sky130_fd_sc_hd__mux2_1
XFILLER_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18058_ _01757_ _01758_ _01759_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__nand3_1
XFILLER_172_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17009_ _09499_ _09506_ _09648_ vssd1 vssd1 vccd1 vccd1 _09649_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20020_ _04891_ _04887_ _04886_ _04890_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__or4b_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20922_ clknet_leaf_18_i_clk _00691_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20853_ clknet_leaf_45_i_clk _00622_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20784_ clknet_leaf_27_i_clk _00553_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_148_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21405_ net326 _01174_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21336_ net257 _01105_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[43\] sky130_fd_sc_hd__dfxtp_1
X_20332__343 clknet_1_1__leaf__03315_ vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__inv_2
XFILLER_190_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21267_ clknet_leaf_89_i_clk _01036_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11020_ rbzero.tex_b0\[48\] rbzero.tex_b0\[47\] _03854_ vssd1 vssd1 vccd1 vccd1 _03859_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21198_ clknet_leaf_4_i_clk _00967_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.mosi_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20149_ clknet_1_1__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__buf_1
XFILLER_106_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20057__95 clknet_1_1__leaf__03045_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__inv_2
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _05591_ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__nand2_1
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _05741_ _07402_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__nand2_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11922_ _04692_ _04694_ _04697_ _04332_ _04371_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__a221o_1
X_15690_ _08054_ vssd1 vssd1 vccd1 vccd1 _08335_ sky130_fd_sc_hd__clkbuf_4
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _05793_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__buf_2
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ rbzero.tex_g1\[15\] _04327_ _04328_ _04265_ vssd1 vssd1 vccd1 vccd1 _04630_
+ sky130_fd_sc_hd__a31o_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _09243_ _08821_ _09028_ _09164_ vssd1 vssd1 vccd1 vccd1 _09927_ sky130_fd_sc_hd__or4_1
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10804_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _03740_ vssd1 vssd1 vccd1 vccd1 _03746_
+ sky130_fd_sc_hd__mux2_1
XFILLER_202_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11784_ rbzero.tex_g0\[59\] rbzero.tex_g0\[58\] _04212_ vssd1 vssd1 vccd1 vccd1 _04562_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14572_ _07095_ _07096_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__nand2_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16311_ _08617_ _08672_ vssd1 vssd1 vccd1 vccd1 _08956_ sky130_fd_sc_hd__nand2_1
XFILLER_185_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13523_ _05991_ _06080_ _06134_ _05978_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__o22a_1
XFILLER_186_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10735_ _03709_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17291_ _04016_ vssd1 vssd1 vccd1 vccd1 _09863_ sky130_fd_sc_hd__buf_4
XFILLER_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19030_ _02646_ vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_185_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16242_ _08885_ _08886_ vssd1 vssd1 vccd1 vccd1 _08887_ sky130_fd_sc_hd__and2_1
XFILLER_146_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10666_ _03673_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__clkbuf_1
X_13454_ _06069_ _06074_ _06089_ _06190_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__a31oi_2
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12405_ _04989_ gpout0.vpos\[5\] _04891_ _04890_ _05143_ net34 vssd1 vssd1 vccd1
+ vccd1 _05172_ sky130_fd_sc_hd__mux4_1
X_16173_ _08816_ _08075_ _08817_ _08784_ vssd1 vssd1 vccd1 vccd1 _08818_ sky130_fd_sc_hd__nor4_1
X_13385_ _06094_ _06096_ _06095_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__a21boi_1
XFILLER_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10597_ rbzero.tex_g1\[56\] rbzero.tex_g1\[57\] _03635_ vssd1 vssd1 vccd1 vccd1 _03637_
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15124_ rbzero.wall_tracer.rayAddendX\[2\] _07781_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07782_ sky130_fd_sc_hd__mux2_1
X_12336_ _04867_ _05081_ net47 vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__a21oi_1
XFILLER_138_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12267_ _04883_ _04884_ _05021_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__mux2_1
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19932_ rbzero.debug_overlay.playerY\[3\] _03223_ vssd1 vssd1 vccd1 vccd1 _03227_
+ sky130_fd_sc_hd__nor2_1
X_15055_ _04029_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__buf_4
X_11218_ gpout0.hpos\[4\] gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__and2_1
XFILLER_141_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14006_ _06659_ _06741_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__nand2_1
X_19863_ _03911_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__buf_4
X_12198_ _04966_ net61 _04967_ net18 vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__o211a_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11149_ rbzero.debug_overlay.playerY\[2\] _03934_ _03935_ rbzero.debug_overlay.playerY\[4\]
+ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a221o_1
X_18814_ _02492_ _02493_ _02487_ _02489_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__o211a_1
X_19794_ rbzero.pov.spi_buffer\[70\] rbzero.pov.spi_buffer\[71\] _03047_ vssd1 vssd1
+ vccd1 vccd1 _03126_ sky130_fd_sc_hd__mux2_1
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18745_ _02434_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__clkbuf_1
X_15957_ _08562_ _08558_ vssd1 vssd1 vccd1 vccd1 _08602_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_1_1__f__03294_ clknet_0__03294_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03294_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14908_ _07591_ _07612_ _07613_ _04039_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__o211a_1
X_18676_ _02369_ _02371_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__xnor2_1
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _08514_ _08530_ vssd1 vssd1 vccd1 vccd1 _08533_ sky130_fd_sc_hd__nor2_1
XFILLER_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17627_ _10085_ _10187_ _10191_ vssd1 vssd1 vccd1 vccd1 _10192_ sky130_fd_sc_hd__a21oi_1
XFILLER_93_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14839_ _07459_ _07444_ _07468_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__o21bai_4
XFILLER_64_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17558_ _09994_ _10002_ _10123_ vssd1 vssd1 vccd1 vccd1 _10124_ sky130_fd_sc_hd__a21bo_1
XFILLER_205_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16509_ _09113_ _09152_ vssd1 vssd1 vccd1 vccd1 _09153_ sky130_fd_sc_hd__xnor2_2
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17489_ _10053_ _10054_ vssd1 vssd1 vccd1 vccd1 _10055_ sky130_fd_sc_hd__nand2_1
XFILLER_177_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19228_ rbzero.spi_registers.vshift\[0\] _02762_ _02764_ _02765_ vssd1 vssd1 vccd1
+ vccd1 _00758_ sky130_fd_sc_hd__o211a_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19159_ rbzero.spi_registers.new_other\[1\] _02712_ vssd1 vssd1 vccd1 vccd1 _02720_
+ sky130_fd_sc_hd__or2_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21121_ net211 _00890_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21052_ clknet_leaf_73_i_clk _00821_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20003_ rbzero.pov.ready_buffer\[7\] _03246_ _03248_ rbzero.debug_overlay.vplaneY\[-2\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__a221o_1
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20905_ clknet_leaf_88_i_clk _00674_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20836_ clknet_opt_10_1_i_clk _00605_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20767_ clknet_leaf_29_i_clk _00536_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10520_ _03596_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_156_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20698_ clknet_leaf_56_i_clk _00482_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _03560_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_148_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13170_ _05800_ _05906_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__or2_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10382_ rbzero.tex_r1\[28\] rbzero.tex_r1\[29\] _03516_ vssd1 vssd1 vccd1 vccd1 _03522_
+ sky130_fd_sc_hd__mux2_1
XFILLER_163_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12121_ _04890_ _04891_ _04892_ gpout0.vpos\[0\] _04852_ _04846_ vssd1 vssd1 vccd1
+ vccd1 _04893_ sky130_fd_sc_hd__mux4_1
X_21319_ net240 _01088_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12052_ rbzero.row_render.texu\[5\] rbzero.row_render.texu\[4\] _03473_ vssd1 vssd1
+ vccd1 vccd1 _04826_ sky130_fd_sc_hd__mux2_1
XFILLER_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11003_ rbzero.tex_b0\[56\] rbzero.tex_b0\[55\] _03843_ vssd1 vssd1 vccd1 vccd1 _03850_
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16860_ _09096_ _08427_ vssd1 vssd1 vccd1 vccd1 _09501_ sky130_fd_sc_hd__nor2_1
XFILLER_89_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15811_ _08442_ _08455_ vssd1 vssd1 vccd1 vccd1 _08456_ sky130_fd_sc_hd__xor2_1
X_16791_ _09085_ _09431_ _09432_ _08235_ vssd1 vssd1 vccd1 vccd1 _09433_ sky130_fd_sc_hd__o31ai_4
XFILLER_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18530_ _02226_ _02227_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__or2_1
X_15742_ _07996_ _08194_ vssd1 vssd1 vccd1 vccd1 _08387_ sky130_fd_sc_hd__nor2_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _05690_ _05634_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__or2_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18461_ _02144_ _02158_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__xnor2_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _04678_ _04679_ _04680_ _04345_ _04253_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__o221a_1
XFILLER_93_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15673_ _08263_ _08264_ _08307_ vssd1 vssd1 vccd1 vccd1 _08318_ sky130_fd_sc_hd__a21o_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12885_ _04001_ _05490_ _05620_ _05621_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__o2bb2a_2
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _09694_ _09701_ _09978_ vssd1 vssd1 vccd1 vccd1 _09979_ sky130_fd_sc_hd__a21bo_1
XFILLER_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _05893_ _07360_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__and2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _04611_ _04612_ _04304_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__mux2_1
X_18392_ _02089_ _02090_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__xor2_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _08331_ _09621_ vssd1 vssd1 vccd1 vccd1 _09910_ sky130_fd_sc_hd__nand2_1
XFILLER_198_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14555_ _07287_ _07288_ _07291_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__o21a_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _04543_ _04544_ _04138_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__mux2_1
XFILLER_201_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20339__349 clknet_1_1__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__inv_2
XFILLER_14_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13506_ _06241_ _06242_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__nand2_1
XFILLER_186_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10718_ _03700_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__clkbuf_1
X_17274_ _09838_ _09840_ _09839_ vssd1 vssd1 vccd1 vccd1 _09848_ sky130_fd_sc_hd__o21bai_2
XFILLER_174_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14486_ _06689_ _06708_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__nor2_1
X_11698_ rbzero.debug_overlay.vplaneY\[-6\] _04475_ _04454_ rbzero.debug_overlay.vplaneY\[-5\]
+ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a221o_1
X_19013_ _02637_ vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__clkbuf_1
X_16225_ _08868_ _08869_ vssd1 vssd1 vccd1 vccd1 _08870_ sky130_fd_sc_hd__or2_1
X_13437_ _05943_ _06000_ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__and2b_1
X_10649_ _03664_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16156_ _08766_ _08800_ vssd1 vssd1 vccd1 vccd1 _08801_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_41_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13368_ _06103_ _06104_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__nand2_1
XFILLER_115_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15107_ _07764_ _07765_ vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__or2_1
X_12319_ _05083_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__clkbuf_4
X_16087_ _08728_ _08731_ vssd1 vssd1 vccd1 vccd1 _08732_ sky130_fd_sc_hd__or2b_1
X_13299_ _06032_ _06033_ _06034_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__nand3_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15038_ _07700_ _07701_ _03914_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__a21oi_1
X_19915_ rbzero.pov.ready_buffer\[52\] _03164_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__nor2_1
XFILLER_190_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_56_i_clk clknet_3_6_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19846_ _03139_ _03160_ _03161_ _03157_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__o211a_1
XFILLER_96_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16989_ _08075_ _08821_ _09028_ _08425_ vssd1 vssd1 vccd1 vccd1 _09629_ sky130_fd_sc_hd__or4_1
XFILLER_7_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19777_ _03117_ vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20084__119 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__inv_2
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18728_ rbzero.wall_tracer.trackDistY\[-9\] _02419_ _02399_ vssd1 vssd1 vccd1 vccd1
+ _02420_ sky130_fd_sc_hd__mux2_1
XFILLER_83_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18659_ _01860_ _09027_ _09350_ _01498_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__o22ai_1
XFILLER_52_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20621_ clknet_leaf_16_i_clk _00405_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.i_row\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_178_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20552_ _03436_ _03439_ _03440_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__a21oi_1
XFILLER_149_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20483_ rbzero.traced_texa\[0\] rbzero.texV\[0\] vssd1 vssd1 vccd1 vccd1 _03383_
+ sky130_fd_sc_hd__or2_1
XFILLER_193_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_7_0_i_clk clknet_2_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_69_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21104_ net194 _00873_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21035_ clknet_leaf_6_i_clk _00804_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready sky130_fd_sc_hd__dfxtp_1
XFILLER_99_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12670_ _05416_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nand2_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _04230_ _04395_ _04399_ _04371_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a211o_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20819_ clknet_leaf_49_i_clk _00588_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_179_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14340_ _07075_ _07076_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__and2_1
XFILLER_168_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11552_ rbzero.tex_r1\[13\] rbzero.tex_r1\[12\] _04291_ vssd1 vssd1 vccd1 vccd1 _04331_
+ sky130_fd_sc_hd__mux2_1
XFILLER_196_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10503_ _03587_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11483_ _04262_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__clkbuf_8
X_14271_ _06245_ _06663_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__nor2_1
XFILLER_11_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ _08637_ _08629_ vssd1 vssd1 vccd1 vccd1 _08655_ sky130_fd_sc_hd__or2b_1
Xclkbuf_1_0__f__03297_ clknet_0__03297_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03297_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10434_ _03482_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__clkbuf_4
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13222_ _05931_ _05911_ _05958_ _05928_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__o211a_1
XFILLER_87_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10365_ rbzero.tex_r1\[36\] rbzero.tex_r1\[37\] _03505_ vssd1 vssd1 vccd1 vccd1 _03513_
+ sky130_fd_sc_hd__mux2_1
XFILLER_151_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13153_ _05773_ _05733_ _05792_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__mux2_1
X_12104_ net4 _04875_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__or2_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17961_ _01560_ _01663_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__xor2_1
XFILLER_151_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13084_ _05815_ _05819_ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__mux2_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12035_ gpout0.hpos\[3\] vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__clkbuf_4
X_16912_ _09117_ _09552_ vssd1 vssd1 vccd1 vccd1 _09553_ sky130_fd_sc_hd__nor2_2
X_19700_ rbzero.pov.spi_buffer\[25\] rbzero.pov.spi_buffer\[26\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03077_ sky130_fd_sc_hd__mux2_1
X_17892_ _08202_ _01475_ _01476_ _08259_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__o22ai_1
Xclkbuf_0__03300_ _03300_ vssd1 vssd1 vccd1 vccd1 clknet_0__03300_ sky130_fd_sc_hd__clkbuf_16
XFILLER_93_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16843_ _09483_ vssd1 vssd1 vccd1 vccd1 _09484_ sky130_fd_sc_hd__clkbuf_4
XFILLER_120_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19562_ rbzero.pov.spi_counter\[3\] rbzero.pov.spi_counter\[2\] _03022_ rbzero.pov.spi_counter\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__a31o_1
X_16774_ _08242_ _09129_ vssd1 vssd1 vccd1 vccd1 _09416_ sky130_fd_sc_hd__and2_1
XFILLER_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13986_ _06720_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__or2b_1
XFILLER_206_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18513_ _02205_ _02206_ _02210_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a21oi_1
X_15725_ _08349_ _08369_ vssd1 vssd1 vccd1 vccd1 _08370_ sky130_fd_sc_hd__xnor2_2
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19493_ _02972_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__clkbuf_1
X_12937_ _05667_ _05650_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__xor2_1
XFILLER_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ _02049_ _02051_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__nor2_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15656_ _07601_ _08148_ _05198_ _08199_ vssd1 vssd1 vccd1 vccd1 _08301_ sky130_fd_sc_hd__and4_1
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12868_ _05563_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__nand2_1
XFILLER_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _07218_ _07323_ _07216_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__a21oi_1
X_18375_ _10094_ _09215_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__nor2_1
X_11819_ rbzero.tex_g1\[51\] rbzero.tex_g1\[50\] _04212_ vssd1 vssd1 vccd1 vccd1 _04596_
+ sky130_fd_sc_hd__mux2_1
X_15587_ _07568_ vssd1 vssd1 vccd1 vccd1 _08232_ sky130_fd_sc_hd__inv_2
XFILLER_15_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ rbzero.wall_tracer.mapY\[7\] _05397_ _05540_ vssd1 vssd1 vccd1 vccd1 _05541_
+ sky130_fd_sc_hd__o21a_1
X_17326_ _09889_ _09893_ _09894_ _09780_ vssd1 vssd1 vccd1 vccd1 _09895_ sky130_fd_sc_hd__a31o_1
XFILLER_186_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14538_ _07233_ _07249_ _07247_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__a21oi_1
XFILLER_159_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257_ _09830_ _09831_ _09832_ vssd1 vssd1 vccd1 vccd1 _09833_ sky130_fd_sc_hd__and3_1
X_14469_ _07131_ _07205_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__nor2_1
X_16208_ _08847_ _08852_ vssd1 vssd1 vccd1 vccd1 _08853_ sky130_fd_sc_hd__nand2_1
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17188_ _09773_ vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16139_ _08519_ _08674_ _08112_ _08377_ vssd1 vssd1 vccd1 vccd1 _08784_ sky130_fd_sc_hd__o22a_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19829_ _03139_ _03147_ _03149_ _02765_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__o211a_1
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21653_ clknet_leaf_37_i_clk _01422_ vssd1 vssd1 vccd1 vccd1 gpout1.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20604_ _03466_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__clkbuf_1
X_21584_ net505 _01353_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20535_ rbzero.traced_texa\[7\] rbzero.texV\[7\] _03422_ vssd1 vssd1 vccd1 vccd1
+ _03427_ sky130_fd_sc_hd__a21o_1
XFILLER_165_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xtop_ew_algofoogle_78 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_78/HI o_rgb[8] sky130_fd_sc_hd__conb_1
Xtop_ew_algofoogle_89 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_89/HI o_rgb[21] sky130_fd_sc_hd__conb_1
XFILLER_137_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20466_ _03362_ _03364_ _03363_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__o21bai_1
XFILLER_192_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21018_ clknet_leaf_9_i_clk _00787_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13840_ _05752_ _05921_ _06053_ _05974_ _05989_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__a32o_1
XFILLER_207_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13771_ _06471_ _06472_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__nand2_1
X_10983_ _03839_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15510_ _08043_ _08055_ vssd1 vssd1 vccd1 vccd1 _08155_ sky130_fd_sc_hd__and2b_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12722_ _05423_ _05428_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__or2_1
X_16490_ _07598_ _08230_ _08147_ _08984_ vssd1 vssd1 vccd1 vccd1 _09134_ sky130_fd_sc_hd__or4_1
XFILLER_128_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15441_ _08076_ _08085_ vssd1 vssd1 vccd1 vccd1 _08086_ sky130_fd_sc_hd__or2_1
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _05403_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18160_ _01860_ _10238_ _09973_ _01737_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__o22ai_1
XFILLER_169_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11604_ _04210_ _04377_ _04382_ _04232_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__a211o_1
X_15372_ _07933_ _07524_ _08016_ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__o21ai_1
XFILLER_12_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12584_ _05297_ _05337_ _05296_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__a21bo_1
XFILLER_196_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17111_ _03555_ _04037_ vssd1 vssd1 vccd1 vccd1 _09749_ sky130_fd_sc_hd__nor2_1
X_14323_ _05982_ _06658_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__nor2_1
XFILLER_157_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11535_ gpout0.vpos\[5\] gpout0.vpos\[4\] vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__or2b_4
X_18091_ rbzero.wall_tracer.trackDistX\[5\] rbzero.wall_tracer.stepDistX\[5\] vssd1
+ vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__or2_1
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17042_ _09409_ _09543_ _09681_ vssd1 vssd1 vccd1 vccd1 _09682_ sky130_fd_sc_hd__a21bo_2
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14254_ _06951_ _06988_ _06990_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__a21o_1
X_11466_ rbzero.tex_r0\[47\] rbzero.tex_r0\[46\] _04213_ vssd1 vssd1 vccd1 vccd1 _04246_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13205_ _05941_ _05910_ _05923_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__o21ai_1
XFILLER_174_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10417_ _03540_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_178_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11397_ gpout0.hpos\[9\] _04158_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__o21a_1
X_14185_ _06666_ _06690_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__nor2_1
XFILLER_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20115__148 clknet_1_1__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__inv_2
XFILLER_152_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13136_ _05791_ _05795_ _05591_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__or3b_1
X_10348_ rbzero.tex_r1\[44\] rbzero.tex_r1\[45\] _03494_ vssd1 vssd1 vccd1 vccd1 _03504_
+ sky130_fd_sc_hd__mux2_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ _02594_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__buf_4
XFILLER_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ _01643_ _01644_ _01646_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__nand3_2
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _05591_ _05803_ _05791_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__mux2_1
XFILLER_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12018_ rbzero.tex_b1\[47\] _04327_ _04328_ _04265_ vssd1 vssd1 vccd1 vccd1 _04793_
+ sky130_fd_sc_hd__a31o_1
X_17875_ _09249_ _01576_ _01577_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__o21ba_1
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16826_ _09082_ _09467_ vssd1 vssd1 vccd1 vccd1 _09468_ sky130_fd_sc_hd__nor2_1
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16757_ _09397_ _09398_ vssd1 vssd1 vccd1 vccd1 _09399_ sky130_fd_sc_hd__xnor2_1
X_19545_ rbzero.pov.sclk_buffer\[2\] rbzero.pov.sclk_buffer\[1\] vssd1 vssd1 vccd1
+ vccd1 _03019_ sky130_fd_sc_hd__nor2b_2
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13969_ _06613_ _06563_ _06600_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__or3_1
XFILLER_74_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15708_ _08022_ _08035_ _08046_ _08112_ vssd1 vssd1 vccd1 vccd1 _08353_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03045_ clknet_0__03045_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03045_
+ sky130_fd_sc_hd__clkbuf_16
X_16688_ _09207_ _09330_ vssd1 vssd1 vccd1 vccd1 _09331_ sky130_fd_sc_hd__xnor2_4
X_19476_ _02938_ _02956_ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__xor2_1
XFILLER_94_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18427_ _02122_ _02124_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__nand2_1
X_15639_ _07924_ vssd1 vssd1 vccd1 vccd1 _08284_ sky130_fd_sc_hd__buf_6
XFILLER_179_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18358_ _01977_ _01997_ _01975_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17309_ _09879_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__clkbuf_1
X_18289_ _08802_ _10139_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__nor2_1
XFILLER_175_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_12_0_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_12_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_200_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21636_ clknet_leaf_41_i_clk _01405_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21567_ net488 _01336_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_166_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11320_ _04069_ _04097_ _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__o21a_1
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20518_ _03411_ _03412_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__nand2_1
X_21498_ net419 _01267_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11251_ rbzero.vga_sync.vsync _03555_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nor2_8
XFILLER_10_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20449_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] _03354_ vssd1 vssd1 vccd1 vccd1
+ _03355_ sky130_fd_sc_hd__o21ai_1
XFILLER_134_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ rbzero.map_rom.f3 rbzero.map_rom.f2 rbzero.map_rom.a6 rbzero.map_rom.i_row\[4\]
+ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__a22o_1
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15990_ _07958_ _08041_ vssd1 vssd1 vccd1 vccd1 _08635_ sky130_fd_sc_hd__or2_1
X_14941_ rbzero.wall_tracer.visualWallDist\[5\] _07618_ vssd1 vssd1 vccd1 vccd1 _07637_
+ sky130_fd_sc_hd__or2_1
XFILLER_102_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17660_ _10215_ _10224_ vssd1 vssd1 vccd1 vccd1 _10225_ sky130_fd_sc_hd__xnor2_1
XFILLER_169_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14872_ rbzero.wall_tracer.stepDistY\[10\] _07586_ _05188_ vssd1 vssd1 vccd1 vccd1
+ _07587_ sky130_fd_sc_hd__mux2_1
X_16611_ _09252_ _09253_ vssd1 vssd1 vccd1 vccd1 _09254_ sky130_fd_sc_hd__nand2_1
X_13823_ _06378_ _06558_ _06559_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__a21o_2
X_17591_ _10011_ _10013_ vssd1 vssd1 vccd1 vccd1 _10157_ sky130_fd_sc_hd__or2b_1
XFILLER_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16542_ _09183_ _09185_ vssd1 vssd1 vccd1 vccd1 _09186_ sky130_fd_sc_hd__xnor2_4
X_19330_ _02821_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__clkbuf_4
X_13754_ _06483_ _06485_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__nand2_1
XFILLER_16_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10966_ rbzero.tex_b1\[9\] rbzero.tex_b1\[10\] _03828_ vssd1 vssd1 vccd1 vccd1 _03831_
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _05451_ _05452_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__nand2_1
X_19261_ _02784_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__clkbuf_1
X_16473_ _08194_ vssd1 vssd1 vccd1 vccd1 _09117_ sky130_fd_sc_hd__buf_4
XFILLER_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13685_ _06379_ _06421_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__nor2_1
X_10897_ _03794_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__clkbuf_1
X_18212_ _01909_ _01910_ _01911_ _05204_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__o31a_1
XFILLER_19_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15424_ rbzero.debug_overlay.playerY\[-3\] _07952_ vssd1 vssd1 vccd1 vccd1 _08069_
+ sky130_fd_sc_hd__nand2_1
X_19192_ rbzero.spi_registers.new_sky\[0\] rbzero.spi_registers.got_new_sky _02711_
+ _02741_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a31o_1
X_12636_ rbzero.map_rom.a6 _05374_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__or2_1
XFILLER_129_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18143_ _10239_ _08423_ _01843_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__or3_1
X_15355_ rbzero.debug_overlay.playerX\[-7\] vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__inv_2
XFILLER_89_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12567_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[9\] vssd1
+ vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__or2_1
XFILLER_102_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14306_ _07042_ _06995_ _07039_ _07038_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__a31o_1
X_18074_ _01773_ _01774_ _01733_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a21oi_1
X_11518_ _04294_ _04297_ _04210_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__mux2_1
XFILLER_117_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15286_ _07929_ _07930_ vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__or2_2
X_12498_ _05251_ rbzero.wall_tracer.trackDistX\[-2\] _05252_ rbzero.wall_tracer.trackDistX\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__o22a_1
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17025_ _09661_ _08047_ _09662_ _09664_ vssd1 vssd1 vccd1 vccd1 _09665_ sky130_fd_sc_hd__or4bb_2
X_14237_ _06844_ _06973_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__and2_1
XFILLER_125_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11449_ _04123_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__buf_4
XFILLER_153_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14168_ _06903_ _06904_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__and2b_1
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _05852_ _05853_ _05855_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a21o_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _06823_ _06834_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__or2b_1
X_18976_ _02618_ vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__clkbuf_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _01622_ _01629_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__xnor2_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17858_ _01457_ _01490_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__nand2_1
XFILLER_187_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16809_ _09347_ _09450_ vssd1 vssd1 vccd1 vccd1 _09451_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17789_ _10247_ _10250_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__nor2_1
XFILLER_82_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19528_ _03003_ _03004_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__nor2_1
XFILLER_207_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19459_ _02927_ _02938_ _02939_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__nor3_1
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21421_ net342 _01190_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21352_ net273 _01121_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21283_ clknet_leaf_37_i_clk _01052_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_2_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20250__269 clknet_1_1__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__inv_2
XFILLER_104_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _03754_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__clkbuf_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ clknet_leaf_3_i_clk _00767_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20144__174 clknet_1_0__leaf__03296_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__inv_2
XFILLER_164_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10751_ _03717_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__clkbuf_4
XFILLER_38_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13470_ _06200_ _06206_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10682_ rbzero.tex_g1\[16\] rbzero.tex_g1\[17\] _03680_ vssd1 vssd1 vccd1 vccd1 _03682_
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ rbzero.hsync vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__inv_2
XFILLER_185_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21619_ clknet_leaf_73_i_clk _01388_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15140_ _07756_ _07789_ _07790_ _07796_ vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__a31o_1
X_12352_ _04154_ _03477_ _05087_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__mux2_1
XFILLER_154_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11303_ _04079_ _04078_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__nand2_1
X_15071_ _07729_ _07731_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__nand2_1
X_12283_ _04867_ _05027_ _05042_ _05049_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__and4_1
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14022_ _06641_ _06642_ _06615_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__a21o_2
XFILLER_88_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11234_ _04018_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__buf_4
XFILLER_136_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18830_ rbzero.wall_tracer.trackDistY\[4\] _02508_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02509_ sky130_fd_sc_hd__mux2_1
XFILLER_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ _03939_ _03952_ _03953_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__o21a_1
XFILLER_136_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18761_ rbzero.wall_tracer.trackDistY\[-5\] _02448_ _02441_ vssd1 vssd1 vccd1 vccd1
+ _02449_ sky130_fd_sc_hd__mux2_1
XFILLER_95_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11096_ rbzero.tex_b0\[12\] rbzero.tex_b0\[11\] _03898_ vssd1 vssd1 vccd1 vccd1 _03899_
+ sky130_fd_sc_hd__mux2_1
X_15973_ _08615_ _08614_ vssd1 vssd1 vccd1 vccd1 _08618_ sky130_fd_sc_hd__and2b_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17712_ _10254_ _10276_ vssd1 vssd1 vccd1 vccd1 _10277_ sky130_fd_sc_hd__xnor2_2
X_14924_ _07621_ _07624_ _07625_ _07620_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__o211a_1
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18692_ _02310_ _02313_ _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__o21a_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17643_ _09249_ _09359_ vssd1 vssd1 vccd1 vccd1 _10208_ sky130_fd_sc_hd__nor2_1
X_14855_ _07433_ _07421_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__nand2_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13806_ _06522_ _06524_ _06526_ _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__or4_1
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17574_ _08872_ _08873_ _09991_ _10139_ vssd1 vssd1 vccd1 vccd1 _10140_ sky130_fd_sc_hd__or4_1
X_14786_ _05884_ _07517_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__nor2_1
XFILLER_205_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11998_ rbzero.tex_b1\[51\] rbzero.tex_b1\[50\] _04250_ vssd1 vssd1 vccd1 vccd1 _04773_
+ sky130_fd_sc_hd__mux2_1
XFILLER_147_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16525_ _08112_ _08329_ _08419_ vssd1 vssd1 vccd1 vccd1 _09169_ sky130_fd_sc_hd__or3_1
X_19313_ rbzero.spi_registers.spi_done _03480_ _02563_ vssd1 vssd1 vccd1 vccd1 _02812_
+ sky130_fd_sc_hd__and3_1
X_13737_ _06473_ _06445_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__xnor2_1
XFILLER_56_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10949_ rbzero.tex_b1\[17\] rbzero.tex_b1\[18\] _03817_ vssd1 vssd1 vccd1 vccd1 _03822_
+ sky130_fd_sc_hd__mux2_1
XFILLER_204_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16456_ _09009_ _09099_ vssd1 vssd1 vccd1 vccd1 _09100_ sky130_fd_sc_hd__xnor2_1
X_19244_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_sky\[0\] _02774_
+ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__mux2_1
X_13668_ _06400_ _06404_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15407_ _07903_ rbzero.wall_tracer.stepDistY\[-10\] vssd1 vssd1 vccd1 vccd1 _08052_
+ sky130_fd_sc_hd__nand2_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19175_ rbzero.spi_registers.got_new_leak _02708_ vssd1 vssd1 vccd1 vccd1 _02731_
+ sky130_fd_sc_hd__and2_1
X_12619_ _05331_ _05335_ _05340_ _05370_ _05372_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__o41ai_4
X_16387_ _08331_ _08420_ vssd1 vssd1 vccd1 vccd1 _09032_ sky130_fd_sc_hd__nand2_1
XFILLER_31_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13599_ _06302_ _06329_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__xnor2_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18126_ _08275_ _09165_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__nor2_1
XFILLER_157_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15338_ _07982_ rbzero.debug_overlay.playerY\[-8\] _05373_ vssd1 vssd1 vccd1 vccd1
+ _07983_ sky130_fd_sc_hd__mux2_1
XFILLER_145_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18057_ _10110_ _09991_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__nor2_1
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15269_ rbzero.debug_overlay.playerX\[-5\] _07898_ vssd1 vssd1 vccd1 vccd1 _07914_
+ sky130_fd_sc_hd__xnor2_2
X_17008_ _09387_ _09390_ _09505_ vssd1 vssd1 vccd1 vccd1 _09648_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18959_ _02609_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__clkbuf_1
X_19605__59 clknet_1_0__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__inv_2
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20921_ clknet_leaf_19_i_clk _00690_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20852_ clknet_leaf_50_i_clk _00621_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20783_ clknet_leaf_72_i_clk _00552_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21404_ net325 _01173_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21335_ net256 _01104_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21266_ clknet_leaf_90_i_clk _01035_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21197_ clknet_leaf_93_i_clk _00966_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12970_ _05593_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__xnor2_1
XFILLER_92_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _04695_ _04696_ _04139_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__mux2_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _07106_ _07107_ _07041_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__and3_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ rbzero.tex_g1\[14\] _04272_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__and2_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _03745_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_207_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14571_ _07306_ _07307_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__nand2_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ rbzero.tex_g0\[56\] _04350_ _04224_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__a21o_1
XFILLER_14_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16310_ _08951_ _08953_ _08954_ vssd1 vssd1 vccd1 vccd1 _08955_ sky130_fd_sc_hd__a21oi_4
XFILLER_14_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13522_ _06080_ _06134_ _05921_ _05989_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__and4bb_1
XFILLER_201_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10734_ rbzero.tex_g0\[56\] rbzero.tex_g0\[55\] _03706_ vssd1 vssd1 vccd1 vccd1 _03709_
+ sky130_fd_sc_hd__mux2_1
X_17290_ _09862_ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_159_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16241_ _08884_ _08865_ _08876_ vssd1 vssd1 vccd1 vccd1 _08886_ sky130_fd_sc_hd__nand3_1
X_13453_ _06077_ _06088_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__and2b_1
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10665_ rbzero.tex_g1\[24\] rbzero.tex_g1\[25\] _03669_ vssd1 vssd1 vccd1 vccd1 _03673_
+ sky130_fd_sc_hd__mux2_1
XFILLER_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12404_ _05141_ _05166_ _05168_ _05170_ _05153_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__o221a_1
XFILLER_167_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16172_ _08674_ _08112_ _08747_ vssd1 vssd1 vccd1 vccd1 _08817_ sky130_fd_sc_hd__nor3_1
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13384_ _06112_ _06118_ _06120_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__a21bo_1
XFILLER_51_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10596_ _03636_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15123_ _07772_ _07773_ _07780_ _07676_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12335_ _05083_ _05082_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__and2b_1
XFILLER_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15054_ _07676_ _07708_ _07709_ _07716_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__a31o_1
X_19931_ rbzero.debug_overlay.playerY\[2\] _03198_ _03226_ _03209_ vssd1 vssd1 vccd1
+ vccd1 _01000_ sky130_fd_sc_hd__o211a_1
XFILLER_99_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12266_ _05032_ _05033_ _05034_ _05024_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__o31a_1
XFILLER_107_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14005_ _06659_ _06741_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__xnor2_1
X_11217_ gpout0.hpos\[5\] vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__clkbuf_4
X_19862_ _03141_ _03171_ _03172_ _03173_ _03155_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__o311a_1
XFILLER_96_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput70 net122 vssd1 vssd1 vccd1 vccd1 o_tex_sclk sky130_fd_sc_hd__clkbuf_1
X_12197_ _04966_ _04666_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__nand2_1
XFILLER_122_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_0_i_clk clknet_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1_0_i_clk sky130_fd_sc_hd__clkbuf_8
X_18813_ _02487_ _02489_ _02492_ _02493_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__a211oi_1
X_11148_ rbzero.debug_overlay.playerY\[2\] _03934_ _03936_ rbzero.debug_overlay.playerX\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19793_ _03125_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18744_ rbzero.wall_tracer.trackDistY\[-7\] _02433_ _02399_ vssd1 vssd1 vccd1 vccd1
+ _02434_ sky130_fd_sc_hd__mux2_1
X_11079_ rbzero.tex_b0\[20\] rbzero.tex_b0\[19\] _03887_ vssd1 vssd1 vccd1 vccd1 _03890_
+ sky130_fd_sc_hd__mux2_1
X_15956_ _08588_ _08600_ vssd1 vssd1 vccd1 vccd1 _08601_ sky130_fd_sc_hd__xor2_2
Xclkbuf_1_1__f__03293_ clknet_0__03293_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03293_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14907_ rbzero.wall_tracer.visualWallDist\[-5\] _07595_ vssd1 vssd1 vccd1 vccd1 _07613_
+ sky130_fd_sc_hd__or2_1
X_18675_ _02259_ _02267_ _02370_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a21oi_1
X_15887_ _08484_ _08479_ vssd1 vssd1 vccd1 vccd1 _08532_ sky130_fd_sc_hd__xnor2_2
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17626_ _10189_ _10190_ vssd1 vssd1 vccd1 vccd1 _10191_ sky130_fd_sc_hd__nand2_1
XFILLER_24_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14838_ _07561_ vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__clkbuf_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17557_ _10001_ _10000_ vssd1 vssd1 vccd1 vccd1 _10123_ sky130_fd_sc_hd__or2b_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14769_ rbzero.wall_tracer.stepDistY\[-9\] _07502_ _07461_ vssd1 vssd1 vccd1 vccd1
+ _07503_ sky130_fd_sc_hd__mux2_1
X_16508_ _09149_ _09151_ vssd1 vssd1 vccd1 vccd1 _09152_ sky130_fd_sc_hd__xnor2_2
X_17488_ _09368_ _09483_ _09910_ vssd1 vssd1 vccd1 vccd1 _10054_ sky130_fd_sc_hd__or3_1
XFILLER_60_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19227_ _02721_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__buf_4
XFILLER_108_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16439_ _09080_ _09082_ _05194_ vssd1 vssd1 vccd1 vccd1 _09084_ sky130_fd_sc_hd__a21o_1
XFILLER_108_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19158_ rbzero.othery\[0\] _02710_ _02719_ _02714_ vssd1 vssd1 vccd1 vccd1 _00734_
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18109_ _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__inv_2
XFILLER_8_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19089_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.mosi _02677_ vssd1
+ vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__mux2_1
XFILLER_133_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21120_ net210 _00889_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21051_ clknet_leaf_71_i_clk _00820_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20002_ rbzero.pov.ready_buffer\[6\] _03239_ _03242_ _04471_ _03254_ vssd1 vssd1
+ vccd1 vccd1 _01043_ sky130_fd_sc_hd__o221a_1
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ clknet_leaf_89_i_clk _00673_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_i_clk clknet_2_1_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20835_ clknet_leaf_66_i_clk _00604_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20766_ clknet_leaf_43_i_clk _00535_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_39_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20697_ clknet_leaf_57_i_clk _00481_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_182_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10450_ rbzero.tex_r0\[63\] rbzero.tex_r0\[62\] _03558_ vssd1 vssd1 vccd1 vccd1 _03560_
+ sky130_fd_sc_hd__mux2_1
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20256__275 clknet_1_0__leaf__03307_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__inv_2
XFILLER_109_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10381_ _03521_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_124_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ gpout0.vpos\[1\] vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__buf_2
XFILLER_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21318_ net239 _01087_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12051_ _04814_ _04824_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__nor2_1
XFILLER_46_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21249_ clknet_leaf_86_i_clk _01018_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_120_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11002_ _03849_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15810_ _08451_ _08453_ _08454_ vssd1 vssd1 vccd1 vccd1 _08455_ sky130_fd_sc_hd__a21oi_1
X_16790_ _07575_ _07579_ _08983_ _07582_ vssd1 vssd1 vccd1 vccd1 _09432_ sky130_fd_sc_hd__o31a_1
XFILLER_19_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15741_ _08384_ _08385_ vssd1 vssd1 vccd1 vccd1 _08386_ sky130_fd_sc_hd__nand2_1
XFILLER_133_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _05632_ _05637_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__or2b_2
XFILLER_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ rbzero.tex_b0\[1\] rbzero.tex_b0\[0\] _04290_ vssd1 vssd1 vccd1 vccd1 _04680_
+ sky130_fd_sc_hd__mux2_1
X_18460_ _02149_ _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__xnor2_1
X_15672_ _08314_ _08315_ _08316_ vssd1 vssd1 vccd1 vccd1 _08317_ sky130_fd_sc_hd__a21bo_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12884_ rbzero.wall_tracer.visualWallDist\[1\] _05571_ _04000_ vssd1 vssd1 vccd1
+ vccd1 _05621_ sky130_fd_sc_hd__a21o_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _08872_ _09977_ _09700_ vssd1 vssd1 vccd1 vccd1 _09978_ sky130_fd_sc_hd__or3_1
XFILLER_61_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14623_ _07358_ _07359_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__xnor2_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ rbzero.tex_g1\[41\] rbzero.tex_g1\[40\] _04350_ vssd1 vssd1 vccd1 vccd1 _04612_
+ sky130_fd_sc_hd__mux2_1
X_18391_ _08257_ _08423_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__nor2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_199_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17342_ _09656_ _09617_ vssd1 vssd1 vccd1 vccd1 _09909_ sky130_fd_sc_hd__or2b_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14554_ _07289_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__nand2_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ rbzero.tex_g0\[23\] rbzero.tex_g0\[22\] _04129_ vssd1 vssd1 vccd1 vccd1 _04544_
+ sky130_fd_sc_hd__mux2_1
XFILLER_159_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13505_ _05974_ _06240_ _06161_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__or3_1
XFILLER_202_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10717_ net47 rbzero.tex_g0\[63\] _03624_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__mux2_1
X_17273_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.stepDistX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _09847_ sky130_fd_sc_hd__nand2_1
XFILLER_147_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14485_ _07172_ _07221_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__xnor2_1
XFILLER_105_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11697_ rbzero.debug_overlay.vplaneY\[-8\] _04466_ _04458_ rbzero.debug_overlay.vplaneY\[-9\]
+ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__a22o_1
XFILLER_174_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16224_ _08170_ _08572_ vssd1 vssd1 vccd1 vccd1 _08869_ sky130_fd_sc_hd__or2_1
X_19012_ rbzero.pov.spi_buffer\[38\] rbzero.pov.ready_buffer\[38\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02637_ sky130_fd_sc_hd__mux2_1
X_13436_ _06082_ _06087_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__nand2_1
X_10648_ rbzero.tex_g1\[32\] rbzero.tex_g1\[33\] _03658_ vssd1 vssd1 vccd1 vccd1 _03664_
+ sky130_fd_sc_hd__mux2_1
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16155_ _08778_ _08798_ _08799_ vssd1 vssd1 vccd1 vccd1 _08800_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13367_ _06100_ _06101_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__xor2_1
XFILLER_182_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10579_ _03627_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _07751_ _07754_ _07763_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__and3_1
X_12318_ _05081_ _05084_ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__and3_1
XFILLER_182_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16086_ _08729_ _08730_ vssd1 vssd1 vccd1 vccd1 _08731_ sky130_fd_sc_hd__xnor2_1
X_13298_ _06032_ _06033_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__a21o_1
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15037_ _07697_ _07698_ _07699_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__o21ai_1
X_19914_ rbzero.debug_overlay.playerY\[-2\] _03198_ _03213_ _03209_ vssd1 vssd1 vccd1
+ vccd1 _00996_ sky130_fd_sc_hd__o211a_1
X_12249_ net18 net19 _05002_ _05009_ _05018_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__o311a_2
XFILLER_64_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19845_ _08067_ _03143_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__nand2_1
XFILLER_96_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19776_ rbzero.pov.spi_buffer\[61\] rbzero.pov.spi_buffer\[62\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03117_ sky130_fd_sc_hd__mux2_1
XFILLER_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16988_ _08821_ _09028_ _08425_ _09243_ vssd1 vssd1 vccd1 vccd1 _09628_ sky130_fd_sc_hd__o22a_1
X_18727_ _09863_ _02417_ _02418_ _09835_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__o31ai_1
X_15939_ _08566_ _08583_ _08492_ vssd1 vssd1 vccd1 vccd1 _08584_ sky130_fd_sc_hd__a21oi_4
XFILLER_37_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18658_ _02263_ _02264_ _02261_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a21boi_1
XFILLER_25_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19595__50 clknet_1_1__leaf__03040_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__inv_2
XFILLER_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17609_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _10175_ sky130_fd_sc_hd__nand2_1
XFILLER_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18589_ _02254_ _02285_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__xor2_1
XFILLER_178_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20620_ clknet_leaf_15_i_clk _00404_ vssd1 vssd1 vccd1 vccd1 rbzero.map_rom.a6 sky130_fd_sc_hd__dfxtp_2
XFILLER_71_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20551_ rbzero.traced_texa\[11\] rbzero.texV\[11\] vssd1 vssd1 vccd1 vccd1 _03440_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_149_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20482_ _03272_ _03381_ _03382_ _03250_ rbzero.texV\[-1\] vssd1 vssd1 vccd1 vccd1
+ _01395_ sky130_fd_sc_hd__a32o_1
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21103_ net193 _00872_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21034_ clknet_leaf_12_i_clk _00803_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_vshift
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _04379_ _04396_ _04397_ _04398_ _04209_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__o221a_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20818_ clknet_leaf_60_i_clk _00587_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-2\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11551_ rbzero.tex_r1\[15\] _04327_ _04328_ _04329_ vssd1 vssd1 vccd1 vccd1 _04330_
+ sky130_fd_sc_hd__a31o_1
X_20749_ clknet_leaf_36_i_clk _00518_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_129_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10502_ rbzero.tex_r0\[38\] rbzero.tex_r0\[37\] _03580_ vssd1 vssd1 vccd1 vccd1 _03587_
+ sky130_fd_sc_hd__mux2_1
XFILLER_156_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14270_ _06762_ _06765_ _06764_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__a21bo_1
XFILLER_52_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11482_ _04211_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__buf_6
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__03296_ clknet_0__03296_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03296_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_155_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13221_ _05688_ _05792_ _05957_ _05778_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a211o_1
X_10433_ _03548_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13152_ _05856_ _05877_ _05888_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__a21o_2
X_10364_ _03512_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_128_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ _04813_ _04811_ _04006_ _03475_ net2 net3 vssd1 vssd1 vccd1 vccd1 _04875_
+ sky130_fd_sc_hd__mux4_1
XFILLER_124_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17960_ _01660_ _01662_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__xnor2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _05797_ _05809_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__nand2_2
XFILLER_152_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16911_ _09551_ vssd1 vssd1 vccd1 vccd1 _09552_ sky130_fd_sc_hd__buf_2
X_12034_ _04808_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_8
X_17891_ _08259_ _08202_ _08157_ _08149_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__or4_1
XFILLER_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16842_ _09482_ vssd1 vssd1 vccd1 vccd1 _09483_ sky130_fd_sc_hd__buf_2
XFILLER_144_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19561_ rbzero.pov.spi_counter\[4\] rbzero.pov.spi_counter\[3\] _03028_ vssd1 vssd1
+ vccd1 vccd1 _03031_ sky130_fd_sc_hd__and3_1
X_16773_ _09407_ _09414_ vssd1 vssd1 vccd1 vccd1 _09415_ sky130_fd_sc_hd__xor2_2
X_13985_ _06719_ _06721_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__and2_1
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18512_ _02208_ _02209_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__nand2_1
XFILLER_20_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15724_ _08367_ _08368_ vssd1 vssd1 vccd1 vccd1 _08369_ sky130_fd_sc_hd__nand2_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ _05657_ _05658_ _05663_ _05672_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__or4_2
XFILLER_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19492_ rbzero.wall_tracer.rayAddendY\[6\] _02971_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _02972_ sky130_fd_sc_hd__mux2_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18443_ _02139_ _02140_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__nor2b_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12867_ rbzero.wall_tracer.visualWallDist\[4\] _05571_ _05572_ vssd1 vssd1 vccd1
+ vccd1 _05604_ sky130_fd_sc_hd__a21o_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ rbzero.wall_tracer.visualWallDist\[-11\] _08148_ _05198_ _08254_ vssd1 vssd1
+ vccd1 vccd1 _08300_ sky130_fd_sc_hd__and4_1
XFILLER_178_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ rbzero.tex_g1\[49\] rbzero.tex_g1\[48\] _04212_ vssd1 vssd1 vccd1 vccd1 _04595_
+ sky130_fd_sc_hd__mux2_1
X_14606_ _07329_ _07330_ _07342_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__nand3b_1
X_18374_ _01939_ _02071_ _02072_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a21o_1
X_15586_ _08230_ rbzero.wall_tracer.stepDistY\[5\] vssd1 vssd1 vccd1 vccd1 _08231_
+ sky130_fd_sc_hd__nand2_1
XFILLER_21_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ rbzero.wall_tracer.mapY\[6\] _05397_ _05538_ vssd1 vssd1 vccd1 vccd1 _05540_
+ sky130_fd_sc_hd__a21bo_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14537_ _07197_ _07195_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__xor2_1
X_17325_ _09890_ _09891_ _09892_ vssd1 vssd1 vccd1 vccd1 _09894_ sky130_fd_sc_hd__o21ai_1
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11749_ rbzero.tex_g0\[9\] rbzero.tex_g0\[8\] _04271_ vssd1 vssd1 vccd1 vccd1 _04527_
+ sky130_fd_sc_hd__mux2_1
XFILLER_144_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14468_ _06724_ _06760_ _07117_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__or3_1
X_17256_ _09823_ _09821_ _09822_ vssd1 vssd1 vccd1 vccd1 _09832_ sky130_fd_sc_hd__a21bo_1
XFILLER_105_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16207_ _08840_ _08846_ vssd1 vssd1 vccd1 vccd1 _08852_ sky130_fd_sc_hd__or2_1
X_13419_ _06154_ _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__or2_1
X_17187_ rbzero.wall_tracer.wall\[1\] rbzero.row_render.wall\[1\] _07830_ vssd1 vssd1
+ vccd1 vccd1 _09773_ sky130_fd_sc_hd__mux2_1
XFILLER_155_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14399_ _06698_ _06740_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__nor2_1
XFILLER_161_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16138_ _08748_ _08745_ _08746_ vssd1 vssd1 vccd1 vccd1 _08783_ sky130_fd_sc_hd__a21oi_1
XFILLER_154_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16069_ _08697_ _08712_ _08713_ vssd1 vssd1 vccd1 vccd1 _08714_ sky130_fd_sc_hd__a21oi_1
XFILLER_115_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19828_ _03148_ _03143_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__nand2_1
XFILLER_25_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19759_ rbzero.pov.spi_buffer\[53\] rbzero.pov.spi_buffer\[54\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03108_ sky130_fd_sc_hd__mux2_1
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21652_ clknet_leaf_37_i_clk _01421_ vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20603_ _02721_ _03464_ _03465_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__and3_1
XFILLER_178_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21583_ net504 _01352_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_123_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20534_ _03424_ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__and2b_1
XFILLER_137_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xtop_ew_algofoogle_79 vssd1 vssd1 vccd1 vccd1 top_ew_algofoogle_79/HI o_rgb[9] sky130_fd_sc_hd__conb_1
XFILLER_193_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20465_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 _03368_
+ sky130_fd_sc_hd__nand2_1
XFILLER_193_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20368__376 clknet_1_1__leaf__03318_ vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__inv_2
XFILLER_88_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21017_ clknet_leaf_3_i_clk _00786_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_other\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20067__104 clknet_1_1__leaf__03289_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__inv_2
XFILLER_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13770_ _06488_ _06506_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__and2_1
X_10982_ rbzero.tex_b1\[1\] rbzero.tex_b1\[2\] _03482_ vssd1 vssd1 vccd1 vccd1 _03839_
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12721_ _05430_ _05433_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__xor2_2
XFILLER_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19574__31 clknet_1_1__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__inv_2
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_i_clk clknet_1_0_1_i_clk vssd1 vssd1 vccd1 vccd1 clknet_2_0_0_i_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15440_ _08084_ _08019_ _08020_ vssd1 vssd1 vccd1 vccd1 _08085_ sky130_fd_sc_hd__or3_2
XFILLER_71_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12652_ _05402_ rbzero.map_rom.i_row\[4\] _05283_ vssd1 vssd1 vccd1 vccd1 _05403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ _04378_ _04380_ _04381_ _04219_ _04230_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__o221a_1
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15371_ _07933_ _08015_ vssd1 vssd1 vccd1 vccd1 _08016_ sky130_fd_sc_hd__nand2_1
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ _05301_ _05336_ _05305_ _05309_ _05299_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__o311ai_4
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_55_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17110_ _03474_ _09748_ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__nor2_1
X_14322_ _07058_ _07001_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__xnor2_1
X_18090_ _09807_ _01790_ _01791_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__or3_2
X_11534_ _04047_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__clkinv_2
XFILLER_172_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17041_ _09114_ _09126_ _09544_ vssd1 vssd1 vccd1 vccd1 _09681_ sky130_fd_sc_hd__or3_1
XFILLER_8_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14253_ _06986_ _06987_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__and2b_1
X_11465_ rbzero.tex_r0\[45\] rbzero.tex_r0\[44\] _04213_ vssd1 vssd1 vccd1 vccd1 _04245_
+ sky130_fd_sc_hd__mux2_1
XFILLER_171_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _05889_ _05900_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__nand2_1
XFILLER_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10416_ rbzero.tex_r1\[12\] rbzero.tex_r1\[13\] _03538_ vssd1 vssd1 vccd1 vccd1 _03540_
+ sky130_fd_sc_hd__mux2_1
XFILLER_178_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14184_ _06919_ _06920_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__nand2_1
XFILLER_174_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11396_ rbzero.row_render.size\[9\] _04155_ rbzero.row_render.size\[10\] vssd1 vssd1
+ vccd1 vccd1 _04176_ sky130_fd_sc_hd__a21oi_1
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13135_ _05705_ _05707_ _05791_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__mux2_1
XFILLER_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10347_ _03503_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_125_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ _02626_ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _10271_ _01645_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nor2_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _05593_ _05706_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__xor2_2
XFILLER_151_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12017_ rbzero.tex_b1\[46\] _04272_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__and2_1
X_17874_ _09391_ _09480_ _09484_ _09249_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__o22a_1
XFILLER_66_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16825_ _09465_ _09466_ vssd1 vssd1 vccd1 vccd1 _09467_ sky130_fd_sc_hd__nor2_1
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19544_ _03914_ _03018_ _03009_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__o21ai_1
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16756_ _08282_ _09103_ vssd1 vssd1 vccd1 vccd1 _09398_ sky130_fd_sc_hd__or2_1
XFILLER_0_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13968_ _06704_ _06658_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__nor2_2
XFILLER_185_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15707_ _08022_ _08034_ _08045_ _08112_ vssd1 vssd1 vccd1 vccd1 _08352_ sky130_fd_sc_hd__or4_1
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03044_ clknet_0__03044_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03044_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_206_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19475_ _02904_ _04471_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__xor2_1
X_12919_ _05650_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__nor2_1
XFILLER_207_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16687_ _09328_ _09329_ vssd1 vssd1 vccd1 vccd1 _09330_ sky130_fd_sc_hd__and2_2
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13899_ _06248_ _06581_ _06583_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__a21o_1
XFILLER_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18426_ _02122_ _02124_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__or2_2
XFILLER_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15638_ _07913_ vssd1 vssd1 vccd1 vccd1 _08283_ sky130_fd_sc_hd__buf_4
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18357_ _02033_ _02055_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15569_ _08002_ _08207_ _08210_ _08213_ _07945_ vssd1 vssd1 vccd1 vccd1 _08214_ sky130_fd_sc_hd__a221o_1
XFILLER_202_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17308_ rbzero.wall_tracer.trackDistX\[-4\] _09878_ _05413_ vssd1 vssd1 vccd1 vccd1
+ _09879_ sky130_fd_sc_hd__mux2_1
X_18288_ _09668_ _09991_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__nor2_1
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17239_ _05413_ vssd1 vssd1 vccd1 vccd1 _09817_ sky130_fd_sc_hd__buf_4
XFILLER_171_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21635_ clknet_leaf_46_i_clk _01404_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21566_ net487 _01335_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_100_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20517_ rbzero.traced_texa\[5\] rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 _03412_
+ sky130_fd_sc_hd__nand2_1
XFILLER_193_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21497_ net418 _01266_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_165_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11250_ rbzero.wall_tracer.state\[0\] vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__inv_2
XFILLER_197_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20448_ rbzero.traced_texa\[-7\] rbzero.texV\[-7\] _03349_ vssd1 vssd1 vccd1 vccd1
+ _03354_ sky130_fd_sc_hd__a21o_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11181_ rbzero.wall_tracer.state\[1\] _03969_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__nand2_1
XFILLER_122_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14940_ rbzero.wall_tracer.trackDistY\[5\] rbzero.wall_tracer.trackDistX\[5\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__mux2_1
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14871_ _07468_ _07585_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__or2b_1
XFILLER_47_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16610_ _08383_ _08111_ _08570_ _08282_ vssd1 vssd1 vccd1 vccd1 _09253_ sky130_fd_sc_hd__o22ai_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13822_ _06278_ _06334_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__xnor2_1
X_17590_ _10088_ _10155_ vssd1 vssd1 vccd1 vccd1 _10156_ sky130_fd_sc_hd__xnor2_1
XFILLER_29_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ _09025_ _09049_ _09184_ vssd1 vssd1 vccd1 vccd1 _09185_ sky130_fd_sc_hd__a21oi_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13753_ _06467_ _06489_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__and2b_1
X_10965_ _03830_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12704_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[11\] vssd1
+ vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__nand2_1
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19260_ rbzero.spi_registers.spi_buffer\[0\] rbzero.spi_registers.new_floor\[0\]
+ _02783_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__mux2_1
XFILLER_91_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16472_ _08962_ _08963_ _09115_ vssd1 vssd1 vccd1 vccd1 _09116_ sky130_fd_sc_hd__a21bo_1
X_13684_ _06391_ _06419_ _06420_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a21oi_2
X_10896_ rbzero.tex_b1\[42\] rbzero.tex_b1\[43\] _03784_ vssd1 vssd1 vccd1 vccd1 _03794_
+ sky130_fd_sc_hd__mux2_1
X_18211_ _01909_ _01910_ _01911_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__o21ai_1
XFILLER_203_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12635_ _05387_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__clkbuf_1
X_15423_ _08066_ _08067_ _05495_ vssd1 vssd1 vccd1 vccd1 _08068_ sky130_fd_sc_hd__mux2_1
X_19191_ _03555_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__buf_6
XFILLER_203_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20121__153 clknet_1_0__leaf__03294_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__inv_2
XFILLER_203_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18142_ _01841_ _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__xnor2_1
X_15354_ _07897_ _07998_ vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__nand2_1
XFILLER_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12566_ rbzero.debug_overlay.facingY\[10\] rbzero.wall_tracer.rayAddendY\[10\] vssd1
+ vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__xor2_1
XFILLER_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11517_ _04295_ _04296_ _04247_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__mux2_1
XFILLER_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14305_ _06882_ _07034_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__nand2_1
XFILLER_102_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18073_ _01733_ _01773_ _01774_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__and3_1
XFILLER_156_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15285_ _05197_ rbzero.wall_tracer.stepDistX\[-4\] vssd1 vssd1 vccd1 vccd1 _07930_
+ sky130_fd_sc_hd__nor2_1
X_12497_ rbzero.wall_tracer.trackDistY\[-3\] vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__inv_2
XFILLER_176_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17024_ _08383_ _09103_ _09663_ vssd1 vssd1 vccd1 vccd1 _09664_ sky130_fd_sc_hd__or3_1
X_14236_ _06964_ _06972_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__xnor2_1
X_11448_ rbzero.tex_r0\[59\] rbzero.tex_r0\[58\] _04214_ vssd1 vssd1 vccd1 vccd1 _04228_
+ sky130_fd_sc_hd__mux2_1
XFILLER_153_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14167_ _06741_ _06888_ _06889_ _06891_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a22o_1
XFILLER_113_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11379_ rbzero.row_render.size\[7\] rbzero.row_render.size\[6\] vssd1 vssd1 vccd1
+ vccd1 _04159_ sky130_fd_sc_hd__xnor2_1
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__clkbuf_4
XFILLER_113_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14098_ _06823_ _06834_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__xnor2_1
X_18975_ rbzero.pov.spi_buffer\[20\] rbzero.pov.ready_buffer\[20\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02618_ sky130_fd_sc_hd__mux2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _01626_ _01628_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__xor2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13049_ _05725_ _05657_ _05658_ _05663_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__or4_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17857_ _10189_ _01452_ _01451_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__o21bai_1
XFILLER_113_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20396__21 clknet_1_1__leaf__03321_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__inv_2
X_16808_ _09448_ _09449_ vssd1 vssd1 vccd1 vccd1 _09450_ sky130_fd_sc_hd__xor2_1
XFILLER_54_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17788_ _01455_ _01491_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__xnor2_1
XFILLER_148_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19527_ _03002_ _03000_ _03001_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__and3_1
X_16739_ _09379_ _09380_ vssd1 vssd1 vccd1 vccd1 _09381_ sky130_fd_sc_hd__nand2_1
XFILLER_207_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20204__228 clknet_1_1__leaf__03302_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__inv_2
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19458_ _02938_ _02939_ _02927_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__o21a_1
XFILLER_90_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18409_ _01936_ _01937_ _01935_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__o21a_2
XFILLER_179_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ _02865_ _02875_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__xnor2_1
X_21420_ net341 _01189_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[63\] sky130_fd_sc_hd__dfxtp_1
X_20096__130 clknet_1_0__leaf__03292_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__inv_2
XFILLER_175_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21351_ net272 _01120_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_108_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21282_ clknet_leaf_38_i_clk _01051_ vssd1 vssd1 vccd1 vccd1 gpout0.vpos\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_162_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20997_ clknet_leaf_11_i_clk _00766_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _03556_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__buf_4
XFILLER_25_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20179__205 clknet_1_0__leaf__03300_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__inv_2
XFILLER_38_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10681_ _03681_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12420_ _05138_ _05140_ _05178_ _05186_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__o2bb2a_2
XFILLER_201_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21618_ clknet_leaf_72_i_clk _01387_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ net28 _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__or2_1
XFILLER_166_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21549_ net470 _01318_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11302_ _04077_ _04080_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__xnor2_1
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15070_ _07730_ rbzero.wall_tracer.rayAddendX\[-1\] vssd1 vssd1 vccd1 vccd1 _07731_
+ sky130_fd_sc_hd__nand2_1
X_12282_ _05042_ _05045_ _05048_ _05050_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a211o_1
XFILLER_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14021_ _06615_ _06641_ _06642_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__nand3_4
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ _03969_ _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__or2_1
XFILLER_134_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11164_ rbzero.wall_tracer.visualWallDist\[11\] vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__clkinv_4
XFILLER_171_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18760_ _09863_ _02446_ _02447_ _09869_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__o31ai_1
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11095_ _03556_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__clkbuf_4
X_15972_ _08550_ _08616_ vssd1 vssd1 vccd1 vccd1 _08617_ sky130_fd_sc_hd__xor2_2
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17711_ _10273_ _10275_ vssd1 vssd1 vccd1 vccd1 _10276_ sky130_fd_sc_hd__xnor2_2
X_14923_ rbzero.wall_tracer.visualWallDist\[-1\] _07618_ vssd1 vssd1 vccd1 vccd1 _07625_
+ sky130_fd_sc_hd__or2_1
X_18691_ _02382_ _02386_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__xor2_4
XFILLER_102_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17642_ _09391_ _10205_ _10206_ vssd1 vssd1 vccd1 vccd1 _10207_ sky130_fd_sc_hd__o21ba_1
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14854_ _07572_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13805_ _05825_ _06031_ _06527_ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__o31a_1
XFILLER_112_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17573_ _10138_ _09565_ _05198_ vssd1 vssd1 vccd1 vccd1 _10139_ sky130_fd_sc_hd__mux2_4
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14785_ _07490_ _07493_ _05952_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__mux2_1
X_11997_ rbzero.tex_b1\[49\] rbzero.tex_b1\[48\] _04250_ vssd1 vssd1 vccd1 vccd1 _04772_
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19312_ rbzero.spi_registers.got_new_other _02730_ _02728_ _02801_ vssd1 vssd1 vccd1
+ vccd1 _00796_ sky130_fd_sc_hd__a31o_1
XFILLER_189_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16524_ _09003_ _09006_ vssd1 vssd1 vccd1 vccd1 _09168_ sky130_fd_sc_hd__nand2_1
XFILLER_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13736_ _06045_ _06016_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__nor2_1
X_10948_ _03821_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19243_ _02773_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__clkbuf_4
X_16455_ _07977_ _08109_ vssd1 vssd1 vccd1 vccd1 _09099_ sky130_fd_sc_hd__nor2_1
X_13667_ _06356_ _06401_ _06402_ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__o22a_1
X_10879_ _03785_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_32_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ rbzero.wall_tracer.side _08049_ _08050_ rbzero.wall_tracer.state\[3\] vssd1
+ vssd1 vccd1 vccd1 _08051_ sky130_fd_sc_hd__o211a_1
X_19174_ rbzero.spi_registers.new_vinf _02726_ _02728_ _02729_ _02730_ vssd1 vssd1
+ vccd1 vccd1 _00739_ sky130_fd_sc_hd__o311a_1
X_12618_ _05327_ _05371_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__nand2_2
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _08416_ _08420_ _08426_ vssd1 vssd1 vccd1 vccd1 _09031_ sky130_fd_sc_hd__a21bo_1
X_13598_ _06278_ _06334_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__nand2_1
XFILLER_12_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18125_ _01824_ _01825_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__xnor2_1
X_12549_ _05301_ _05302_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__nor2_1
X_15337_ rbzero.debug_overlay.playerY\[-8\] rbzero.debug_overlay.playerY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__xor2_1
XFILLER_144_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18056_ _08895_ _08767_ _01524_ _10139_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__or4_1
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _02406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ _07912_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__clkbuf_4
X_17007_ _09639_ _09646_ vssd1 vssd1 vccd1 vccd1 _09647_ sky130_fd_sc_hd__xnor2_1
XFILLER_144_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14219_ _06924_ _06930_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__or2b_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15199_ _07835_ _07838_ _07836_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__a21boi_1
XFILLER_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18958_ rbzero.pov.spi_buffer\[12\] rbzero.pov.ready_buffer\[12\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02609_ sky130_fd_sc_hd__mux2_1
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17909_ _01507_ _01509_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__nor2_1
X_18889_ rbzero.spi_registers.spi_counter\[3\] vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__inv_2
XFILLER_55_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20920_ clknet_leaf_19_i_clk _00689_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20128__159 clknet_1_1__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__inv_2
XFILLER_148_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20851_ clknet_leaf_50_i_clk _00620_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20782_ clknet_leaf_71_i_clk _00551_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21403_ net324 _01172_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21334_ net255 _01103_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_163_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21265_ clknet_leaf_89_i_clk _01034_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20216_ clknet_1_1__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__buf_1
XFILLER_132_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21196_ clknet_leaf_93_i_clk _00965_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11920_ rbzero.tex_b0\[31\] rbzero.tex_b0\[30\] _04271_ vssd1 vssd1 vccd1 vccd1 _04696_
+ sky130_fd_sc_hd__mux2_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _04610_ _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__nor2_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ rbzero.tex_g0\[24\] rbzero.tex_g0\[23\] _03740_ vssd1 vssd1 vccd1 vccd1 _03745_
+ sky130_fd_sc_hd__mux2_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14570_ _07295_ _07300_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__xor2_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11782_ rbzero.tex_g0\[57\] _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__and3_1
XFILLER_54_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20390__16 clknet_1_1__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__inv_2
X_10733_ _03708_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__clkbuf_1
X_13521_ _05990_ _06067_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__or2_1
XFILLER_207_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16240_ _08865_ _08876_ _08884_ vssd1 vssd1 vccd1 vccd1 _08885_ sky130_fd_sc_hd__a21o_1
X_13452_ _06152_ _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__xnor2_1
XFILLER_185_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10664_ _03672_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12403_ _05149_ _05169_ _05145_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a21o_1
XFILLER_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16171_ _08594_ vssd1 vssd1 vccd1 vccd1 _08816_ sky130_fd_sc_hd__clkbuf_4
X_13383_ _06045_ _06114_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__or3_1
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ rbzero.tex_g1\[57\] rbzero.tex_g1\[58\] _03635_ vssd1 vssd1 vccd1 vccd1 _03636_
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12334_ net31 _05099_ _05101_ _04867_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__or4b_1
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15122_ _07778_ _07779_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__xor2_1
XFILLER_86_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15053_ _07676_ _07715_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__nor2_1
X_19930_ rbzero.pov.ready_buffer\[55\] _03141_ _03192_ _03225_ vssd1 vssd1 vccd1 vccd1
+ _03226_ sky130_fd_sc_hd__a211o_1
X_12265_ net24 vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__inv_2
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20233__254 clknet_1_0__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__inv_2
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14004_ _06704_ _06740_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__nor2_1
XFILLER_107_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11216_ _04001_ _04002_ _04003_ _03914_ rbzero.wall_tracer.state\[0\] vssd1 vssd1
+ vccd1 vccd1 _00011_ sky130_fd_sc_hd__a311o_1
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19861_ rbzero.pov.ready_buffer\[69\] _03145_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__or2_1
X_12196_ _04961_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__clkbuf_4
Xoutput60 net60 vssd1 vssd1 vccd1 vccd1 o_reset sky130_fd_sc_hd__buf_2
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 o_vsync sky130_fd_sc_hd__buf_2
XFILLER_122_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18812_ rbzero.wall_tracer.trackDistY\[2\] rbzero.wall_tracer.stepDistY\[2\] vssd1
+ vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__nor2_1
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ rbzero.map_rom.f1 vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__clkinv_2
XFILLER_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19792_ rbzero.pov.spi_buffer\[69\] rbzero.pov.spi_buffer\[70\] _03047_ vssd1 vssd1
+ vccd1 vccd1 _03125_ sky130_fd_sc_hd__mux2_1
XFILLER_96_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18743_ _02431_ _02432_ _09851_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__o21ai_1
XFILLER_114_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03292_ clknet_0__03292_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03292_
+ sky130_fd_sc_hd__clkbuf_16
X_11078_ _03889_ vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__clkbuf_1
X_15955_ _08589_ _08598_ _08599_ vssd1 vssd1 vccd1 vccd1 _08600_ sky130_fd_sc_hd__a21oi_2
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14906_ rbzero.wall_tracer.trackDistY\[-5\] rbzero.wall_tracer.trackDistX\[-5\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__mux2_1
X_18674_ _02265_ _02266_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__and2b_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15886_ _08514_ _08530_ vssd1 vssd1 vccd1 vccd1 _08531_ sky130_fd_sc_hd__xor2_2
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17625_ _10064_ _10067_ _10188_ vssd1 vssd1 vccd1 vccd1 _10190_ sky130_fd_sc_hd__nand3_1
X_14837_ rbzero.wall_tracer.stepDistY\[1\] _07560_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07561_ sky130_fd_sc_hd__mux2_1
XFILLER_63_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17556_ _10112_ _10121_ vssd1 vssd1 vccd1 vccd1 _10122_ sky130_fd_sc_hd__xnor2_2
XFILLER_45_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14768_ _07487_ _07455_ _07488_ _07501_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__a211o_1
XFILLER_108_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_205_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16507_ _08970_ _08994_ _09150_ vssd1 vssd1 vccd1 vccd1 _09151_ sky130_fd_sc_hd__a21bo_1
X_13719_ _06454_ _06439_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__or2b_1
X_17487_ _09368_ _09480_ _09483_ _08329_ vssd1 vssd1 vccd1 vccd1 _10053_ sky130_fd_sc_hd__o22ai_1
XFILLER_177_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14699_ _05892_ _07395_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__nand2_1
XFILLER_60_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19226_ rbzero.spi_registers.new_vshift\[0\] _02763_ vssd1 vssd1 vccd1 vccd1 _02764_
+ sky130_fd_sc_hd__or2_1
XFILLER_177_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16438_ _09080_ _09082_ vssd1 vssd1 vccd1 vccd1 _09083_ sky130_fd_sc_hd__nor2_1
XFILLER_176_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19157_ rbzero.spi_registers.new_other\[0\] _02712_ vssd1 vssd1 vccd1 vccd1 _02719_
+ sky130_fd_sc_hd__or2_1
X_16369_ _08359_ _08360_ vssd1 vssd1 vccd1 vccd1 _09014_ sky130_fd_sc_hd__nand2_1
XFILLER_145_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18108_ _01808_ _01704_ _01702_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__a21oi_1
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19088_ _02676_ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__buf_4
XFILLER_127_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18039_ _01738_ _01740_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__nand2_1
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21050_ clknet_leaf_75_i_clk _00819_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendY\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_193_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20001_ rbzero.pov.ready_buffer\[5\] _03246_ _03248_ rbzero.debug_overlay.vplaneY\[-4\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__a221o_1
XFILLER_87_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20903_ clknet_leaf_88_i_clk _00672_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20834_ clknet_leaf_66_i_clk _00603_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20765_ clknet_leaf_42_i_clk _00534_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20696_ clknet_leaf_57_i_clk _00480_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10380_ rbzero.tex_r1\[29\] rbzero.tex_r1\[30\] _03516_ vssd1 vssd1 vccd1 vccd1 _03521_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21317_ net238 _01086_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12050_ rbzero.row_render.texu\[1\] rbzero.row_render.texu\[0\] _03473_ vssd1 vssd1
+ vccd1 vccd1 _04824_ sky130_fd_sc_hd__mux2_1
X_21248_ clknet_leaf_86_i_clk _01017_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_46_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11001_ rbzero.tex_b0\[57\] rbzero.tex_b0\[56\] _03843_ vssd1 vssd1 vccd1 vccd1 _03849_
+ sky130_fd_sc_hd__mux2_1
XFILLER_117_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21179_ clknet_leaf_7_i_clk _00948_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__04835_ clknet_0__04835_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__04835_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_120_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15740_ _07977_ _08276_ _07981_ _07989_ vssd1 vssd1 vccd1 vccd1 _08385_ sky130_fd_sc_hd__or4_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _05638_ _05649_ _05688_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__or3_1
XFILLER_133_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ rbzero.tex_b0\[2\] _04262_ _04126_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a21o_1
X_15671_ _07913_ _07924_ _07995_ _07932_ vssd1 vssd1 vccd1 vccd1 _08316_ sky130_fd_sc_hd__or4_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12883_ _04030_ _05332_ _05341_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__and3_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _09976_ vssd1 vssd1 vccd1 vccd1 _09977_ sky130_fd_sc_hd__clkbuf_4
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14622_ _07304_ _07308_ _07315_ _07302_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__a31o_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ rbzero.tex_g1\[43\] rbzero.tex_g1\[42\] _04350_ vssd1 vssd1 vccd1 vccd1 _04611_
+ sky130_fd_sc_hd__mux2_1
X_18390_ _02087_ _02088_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__nand2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _09609_ _09612_ _09907_ vssd1 vssd1 vccd1 vccd1 _09908_ sky130_fd_sc_hd__a21o_2
XFILLER_144_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14553_ _07287_ _07288_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__xor2_1
X_11765_ rbzero.tex_g0\[21\] rbzero.tex_g0\[20\] _04129_ vssd1 vssd1 vccd1 vccd1 _04543_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10716_ _03699_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__clkbuf_1
X_13504_ _06239_ _06240_ _06202_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__o21bai_1
XFILLER_186_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17272_ rbzero.wall_tracer.trackDistX\[-7\] rbzero.wall_tracer.stepDistX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _09846_ sky130_fd_sc_hd__or2_1
XFILLER_158_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11696_ _04420_ _04447_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__and2_2
X_14484_ _07176_ _07178_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__xor2_1
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19011_ _02636_ vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__clkbuf_1
X_16223_ _08180_ _08491_ vssd1 vssd1 vccd1 vccd1 _08868_ sky130_fd_sc_hd__or2_1
X_10647_ _03663_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__clkbuf_1
X_13435_ _06170_ _06171_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__xor2_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16154_ _08779_ _08797_ vssd1 vssd1 vccd1 vccd1 _08799_ sky130_fd_sc_hd__nor2_1
X_13366_ _05939_ _06016_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nor2_1
X_10578_ rbzero.tex_r0\[2\] rbzero.tex_r0\[1\] _03624_ vssd1 vssd1 vccd1 vccd1 _03627_
+ sky130_fd_sc_hd__mux2_1
XFILLER_182_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15105_ _07751_ _07754_ _07763_ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__a21oi_1
X_12317_ net29 net28 vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__nor2_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16085_ _08124_ _08490_ _07924_ vssd1 vssd1 vccd1 vccd1 _08730_ sky130_fd_sc_hd__a21oi_1
X_13297_ _05988_ _05980_ _05991_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12248_ _04972_ _05011_ _05017_ net18 vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__a211o_1
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15036_ _07697_ _07698_ _07699_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__or3_1
X_19913_ _08080_ _02823_ _03197_ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__o211ai_1
XFILLER_69_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19844_ rbzero.pov.ready_buffer\[65\] _08066_ _03146_ vssd1 vssd1 vccd1 vccd1 _03160_
+ sky130_fd_sc_hd__mux2_1
XFILLER_110_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12179_ gpout0.vpos\[4\] gpout0.vpos\[5\] _04891_ gpout0.vpos\[9\] net8 net10 vssd1
+ vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__mux4_1
XFILLER_69_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19775_ _03116_ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__clkbuf_1
X_16987_ _08823_ _09164_ vssd1 vssd1 vccd1 vccd1 _09627_ sky130_fd_sc_hd__nor2_1
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18726_ _02414_ _02415_ _02416_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a21oi_1
X_15938_ _08568_ _08582_ vssd1 vssd1 vccd1 vccd1 _08583_ sky130_fd_sc_hd__or2b_1
XFILLER_37_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18657_ _02144_ _02246_ _02352_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__a21oi_1
X_15869_ _08451_ _08453_ vssd1 vssd1 vccd1 vccd1 _08514_ sky130_fd_sc_hd__xnor2_2
XFILLER_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17608_ rbzero.wall_tracer.trackDistX\[1\] rbzero.wall_tracer.stepDistX\[1\] vssd1
+ vssd1 vccd1 vccd1 _10174_ sky130_fd_sc_hd__or2_1
X_18588_ _02268_ _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__xor2_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ _08178_ _09674_ _09965_ _10104_ vssd1 vssd1 vccd1 vccd1 _10105_ sky130_fd_sc_hd__o31a_1
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20550_ _09750_ _03438_ _03439_ _03250_ rbzero.texV\[10\] vssd1 vssd1 vccd1 vccd1
+ _01406_ sky130_fd_sc_hd__a32o_1
XFILLER_177_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19209_ _09753_ _02752_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__and2_1
XFILLER_193_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20481_ _03378_ _03379_ _03373_ _03377_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__a211o_1
XFILLER_193_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21102_ net192 _00871_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[42\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21033_ clknet_leaf_13_i_clk _00802_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20262__280 clknet_1_0__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__inv_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20817_ clknet_leaf_59_i_clk _00586_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-3\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_196_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11550_ _04126_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__buf_4
X_20748_ clknet_leaf_36_i_clk _00517_ vssd1 vssd1 vccd1 vccd1 gpout0.hpos\[0\] sky130_fd_sc_hd__dfxtp_2
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ _03586_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11481_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _04213_ vssd1 vssd1 vccd1 vccd1 _04261_
+ sky130_fd_sc_hd__mux2_1
XFILLER_168_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20679_ clknet_leaf_44_i_clk _00463_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[8\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13220_ _05640_ _05792_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__03295_ clknet_0__03295_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03295_
+ sky130_fd_sc_hd__clkbuf_16
X_10432_ rbzero.tex_r1\[4\] rbzero.tex_r1\[5\] _03538_ vssd1 vssd1 vccd1 vccd1 _03548_
+ sky130_fd_sc_hd__mux2_1
XFILLER_137_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13151_ _05700_ _05879_ _05881_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__a211oi_4
XFILLER_100_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10363_ rbzero.tex_r1\[37\] rbzero.tex_r1\[38\] _03505_ vssd1 vssd1 vccd1 vccd1 _03512_
+ sky130_fd_sc_hd__mux2_1
XFILLER_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12102_ net5 net4 _04873_ net6 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__a31o_1
XFILLER_2_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13082_ _05816_ _05818_ _05806_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__mux2_1
XFILLER_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16910_ _08237_ _09279_ vssd1 vssd1 vccd1 vccd1 _09551_ sky130_fd_sc_hd__and2_1
X_12033_ _04314_ _04807_ _04521_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__o21a_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17890_ _01499_ _01501_ _01497_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__a21bo_1
XFILLER_132_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16841_ _05211_ _09481_ vssd1 vssd1 vccd1 vccd1 _09482_ sky130_fd_sc_hd__or2_1
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19560_ rbzero.pov.spi_counter\[3\] _03028_ _03030_ _03026_ vssd1 vssd1 vccd1 vccd1
+ _00825_ sky130_fd_sc_hd__o211a_1
XFILLER_207_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16772_ _09408_ _09413_ vssd1 vssd1 vccd1 vccd1 _09414_ sky130_fd_sc_hd__xnor2_2
X_20345__355 clknet_1_0__leaf__03316_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__inv_2
XFILLER_207_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13984_ _06710_ _06713_ _06718_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__nand3_1
XFILLER_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18511_ _02078_ _02081_ _02207_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__nand3_1
X_15723_ _08350_ _08351_ _08366_ vssd1 vssd1 vccd1 vccd1 _08368_ sky130_fd_sc_hd__nand3_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19491_ _02967_ _02970_ _04033_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__mux2_1
X_12935_ _05665_ _05666_ _05670_ _05671_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__a22o_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18442_ _10271_ _02028_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__nand2_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _08256_ _08258_ vssd1 vssd1 vccd1 vccd1 _08299_ sky130_fd_sc_hd__xnor2_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12866_ _04031_ _05372_ _05602_ _04001_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__a211o_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14605_ _07340_ _07341_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__and2_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _01498_ _09027_ _09162_ _10239_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__o22a_1
X_11817_ _04594_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_8
XFILLER_57_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _08002_ vssd1 vssd1 vccd1 vccd1 _08230_ sky130_fd_sc_hd__clkbuf_4
XFILLER_30_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12797_ rbzero.wall_tracer.mapY\[7\] _05397_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__and2_1
XFILLER_159_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17324_ _09890_ _09891_ _09892_ vssd1 vssd1 vccd1 vccd1 _09893_ sky130_fd_sc_hd__or3_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _07250_ _07272_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__or2_1
X_11748_ _04523_ _04524_ _04525_ _04139_ _04208_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__o221a_1
XFILLER_187_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17255_ rbzero.wall_tracer.trackDistX\[-9\] rbzero.wall_tracer.stepDistX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _09831_ sky130_fd_sc_hd__nand2_1
XFILLER_175_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14467_ _06689_ _06761_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__or2_1
XFILLER_128_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11679_ _04434_ _04447_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__and2_2
XFILLER_146_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16206_ _08850_ vssd1 vssd1 vccd1 vccd1 _08851_ sky130_fd_sc_hd__inv_2
X_13418_ _06015_ _06031_ _05982_ _05974_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__o22a_1
X_17186_ _09772_ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__clkbuf_1
X_14398_ _07114_ _07127_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__or2_1
XFILLER_154_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16137_ _08748_ _08745_ _08746_ vssd1 vssd1 vccd1 vccd1 _08782_ sky130_fd_sc_hd__and3_1
XFILLER_128_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13349_ _06081_ _06085_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__xnor2_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20090__125 clknet_1_0__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__inv_2
XFILLER_115_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16068_ _08698_ _08711_ vssd1 vssd1 vccd1 vccd1 _08713_ sky130_fd_sc_hd__and2b_1
XFILLER_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15019_ rbzero.debug_overlay.vplaneX\[-7\] rbzero.wall_tracer.rayAddendX\[-7\] vssd1
+ vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__nor2_1
XFILLER_116_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19827_ rbzero.debug_overlay.playerX\[-8\] vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__inv_2
XFILLER_84_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19758_ _03107_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18709_ rbzero.wall_tracer.trackDistY\[-12\] rbzero.wall_tracer.stepDistY\[-12\]
+ _02401_ _02402_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__and4_1
XFILLER_204_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19689_ _03071_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03289_ _03289_ vssd1 vssd1 vccd1 vccd1 clknet_0__03289_ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21651_ clknet_leaf_38_i_clk _01420_ vssd1 vssd1 vccd1 vccd1 gpout0.clk_div\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20602_ gpout2.clk_div\[0\] gpout2.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__or2_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21582_ net503 _01351_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20533_ rbzero.traced_texa\[8\] rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _03425_
+ sky130_fd_sc_hd__nand2_1
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20464_ rbzero.traced_texa\[-3\] rbzero.texV\[-3\] vssd1 vssd1 vccd1 vccd1 _03367_
+ sky130_fd_sc_hd__or2_1
XFILLER_4_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21016_ clknet_leaf_8_i_clk _00785_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.got_new_leak
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10981_ _03838_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12720_ _05421_ _05467_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__xnor2_1
XFILLER_167_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12651_ rbzero.debug_overlay.playerY\[4\] _05401_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05402_ sky130_fd_sc_hd__mux2_1
XFILLER_203_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11602_ rbzero.tex_r1\[59\] rbzero.tex_r1\[58\] _04338_ vssd1 vssd1 vccd1 vccd1 _04381_
+ sky130_fd_sc_hd__mux2_1
XFILLER_130_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12582_ _05289_ _05295_ _05303_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__and3_1
X_15370_ _05351_ _05475_ _07893_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__mux2_1
XFILLER_168_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14321_ _07055_ _07057_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__xnor2_1
X_11533_ _04206_ _04312_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__nand2_1
XFILLER_183_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17040_ _09659_ _09679_ vssd1 vssd1 vccd1 vccd1 _09680_ sky130_fd_sc_hd__xnor2_2
XFILLER_172_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11464_ _04121_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__buf_4
X_14252_ _06951_ _06962_ _06984_ _06988_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__or4_1
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _03539_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__clkbuf_1
X_13203_ _05923_ _05939_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__xnor2_4
X_11395_ _04154_ _04157_ _04158_ gpout0.hpos\[9\] _04174_ vssd1 vssd1 vccd1 vccd1
+ _04175_ sky130_fd_sc_hd__a221o_1
X_14183_ _06709_ _06918_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__or2_1
XFILLER_180_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10346_ rbzero.tex_r1\[45\] rbzero.tex_r1\[46\] _03494_ vssd1 vssd1 vccd1 vccd1 _03503_
+ sky130_fd_sc_hd__mux2_1
X_13134_ _05700_ _05703_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__nor2_2
X_18991_ rbzero.pov.spi_buffer\[28\] rbzero.pov.ready_buffer\[28\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02626_ sky130_fd_sc_hd__mux2_1
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17942_ _10133_ _10135_ _10126_ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__a21boi_2
XFILLER_152_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _05710_ _05715_ _05718_ _05713_ _05777_ _05801_ vssd1 vssd1 vccd1 vccd1 _05802_
+ sky130_fd_sc_hd__mux4_1
XFILLER_124_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12016_ rbzero.tex_b1\[45\] rbzero.tex_b1\[44\] _04392_ vssd1 vssd1 vccd1 vccd1 _04791_
+ sky130_fd_sc_hd__mux2_1
X_17873_ _09391_ _09351_ _09483_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__or3_1
XFILLER_39_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16824_ _09463_ _09464_ vssd1 vssd1 vccd1 vccd1 _09466_ sky130_fd_sc_hd__and2_1
XFILLER_94_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19543_ rbzero.wall_tracer.rayAddendY\[11\] _03017_ vssd1 vssd1 vccd1 vccd1 _03018_
+ sky130_fd_sc_hd__xnor2_1
X_16755_ _09395_ _09396_ vssd1 vssd1 vccd1 vccd1 _09397_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13967_ _06031_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15706_ _08323_ _08317_ vssd1 vssd1 vccd1 vccd1 _08351_ sky130_fd_sc_hd__or2b_1
XFILLER_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_206_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03043_ clknet_0__03043_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03043_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19474_ _07678_ _02953_ _02954_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__and3_1
XFILLER_59_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12918_ _05652_ _05654_ _05567_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a21oi_1
X_16686_ _09208_ _09327_ vssd1 vssd1 vccd1 vccd1 _09329_ sky130_fd_sc_hd__or2_1
X_20404__5 clknet_1_1__leaf__03037_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__inv_2
X_13898_ _06586_ _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__xnor2_2
XFILLER_181_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18425_ _02006_ _02008_ _02123_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__o21a_1
XFILLER_206_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15637_ _07977_ vssd1 vssd1 vccd1 vccd1 _08282_ sky130_fd_sc_hd__clkbuf_4
XFILLER_59_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12849_ _05570_ _05360_ _05585_ _05561_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__o211a_1
XFILLER_181_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18356_ _02035_ _02054_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__xnor2_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15568_ _08002_ _08212_ vssd1 vssd1 vccd1 vccd1 _08213_ sky130_fd_sc_hd__nor2_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17307_ _09812_ _09876_ _09877_ vssd1 vssd1 vccd1 vccd1 _09878_ sky130_fd_sc_hd__o21ai_1
X_14519_ _07231_ _07255_ _05752_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__o21a_1
X_18287_ _01985_ _01986_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__and2_1
XFILLER_175_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15499_ _08138_ _08142_ vssd1 vssd1 vccd1 vccd1 _08144_ sky130_fd_sc_hd__nor2_1
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17238_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.stepDistX\[-12\]
+ _09813_ _09814_ vssd1 vssd1 vccd1 vccd1 _09816_ sky130_fd_sc_hd__a22oi_1
XFILLER_116_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17169_ rbzero.traced_texa\[-2\] _09768_ _09769_ rbzero.wall_tracer.visualWallDist\[-2\]
+ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__a22o_1
XFILLER_155_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21634_ clknet_leaf_46_i_clk _01403_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_139_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21565_ net486 _01334_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20374__381 clknet_1_0__leaf__03319_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__inv_2
X_20516_ rbzero.traced_texa\[5\] rbzero.texV\[5\] vssd1 vssd1 vccd1 vccd1 _03411_
+ sky130_fd_sc_hd__or2_1
X_21496_ net417 _01265_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20447_ _03351_ _03352_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__and2b_1
XFILLER_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11180_ _03955_ _03968_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__and2_1
XFILLER_133_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14870_ _05737_ _05736_ _07584_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__or3_2
XFILLER_76_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13821_ _06425_ _06555_ _06557_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__a21bo_1
XFILLER_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16540_ _09022_ _09024_ vssd1 vssd1 vccd1 vccd1 _09184_ sky130_fd_sc_hd__nor2_1
X_13752_ _06468_ _06482_ _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__a21bo_1
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10964_ rbzero.tex_b1\[10\] rbzero.tex_b1\[11\] _03828_ vssd1 vssd1 vccd1 vccd1 _03830_
+ sky130_fd_sc_hd__mux2_1
X_12703_ rbzero.debug_overlay.facingX\[10\] rbzero.wall_tracer.rayAddendX\[11\] vssd1
+ vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__or2_1
X_16471_ _08282_ _09114_ _08964_ vssd1 vssd1 vccd1 vccd1 _09115_ sky130_fd_sc_hd__or3_1
XFILLER_16_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13683_ _06418_ _06393_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__and2b_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10895_ _03793_ vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__clkbuf_1
X_18210_ _01793_ _01795_ _01794_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__a21boi_1
X_15422_ rbzero.debug_overlay.playerX\[-3\] vssd1 vssd1 vccd1 vccd1 _08067_ sky130_fd_sc_hd__inv_2
XFILLER_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19190_ rbzero.spi_registers.got_new_sky _02707_ vssd1 vssd1 vccd1 vccd1 _02740_
+ sky130_fd_sc_hd__nand2_2
X_12634_ _05386_ _03933_ _05284_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__mux2_1
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18141_ _08257_ _01476_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__nor2_1
XFILLER_145_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15353_ rbzero.debug_overlay.playerX\[-8\] rbzero.debug_overlay.playerX\[-9\] rbzero.debug_overlay.playerX\[-7\]
+ vssd1 vssd1 vccd1 vccd1 _07998_ sky130_fd_sc_hd__o21ai_1
XFILLER_169_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12565_ _05308_ _05312_ _05314_ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__o211a_1
XFILLER_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14304_ _06995_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__xor2_4
X_18072_ _01770_ _01771_ _01772_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a21o_1
X_11516_ rbzero.tex_r0\[23\] rbzero.tex_r0\[22\] _04291_ vssd1 vssd1 vccd1 vccd1 _04296_
+ sky130_fd_sc_hd__mux2_1
XFILLER_89_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15284_ _07925_ _07927_ _07928_ vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__a21oi_1
X_12496_ rbzero.wall_tracer.trackDistY\[-2\] vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__inv_2
XFILLER_171_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17023_ _08202_ _08203_ _08129_ vssd1 vssd1 vccd1 vccd1 _09663_ sky130_fd_sc_hd__a21o_1
XFILLER_172_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14235_ _06938_ _06971_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__and2_1
X_11447_ rbzero.tex_r0\[56\] _04214_ _04226_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__a21o_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11378_ rbzero.row_render.size\[9\] _04155_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__nor2_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14166_ _06853_ _06902_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__or2_1
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10329_ _03482_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__clkbuf_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _05812_ _05821_ _05799_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__mux2_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14097_ _06825_ _06832_ _06833_ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__a21o_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _02617_ vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _09674_ _09417_ _01504_ _01627_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__o31a_1
XFILLER_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13048_ _05701_ _05682_ _05784_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__or3_1
XFILLER_100_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17856_ _01553_ _01559_ rbzero.wall_tracer.trackDistX\[3\] _10036_ vssd1 vssd1 vccd1
+ vccd1 _00592_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16807_ _09239_ _09317_ _09315_ vssd1 vssd1 vccd1 vccd1 _09449_ sky130_fd_sc_hd__a21oi_1
XFILLER_54_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17787_ _01457_ _01490_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__xnor2_1
XFILLER_19_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14999_ rbzero.wall_tracer.stepDistX\[6\] _07571_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07670_ sky130_fd_sc_hd__mux2_1
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16738_ _09263_ _09349_ _09378_ vssd1 vssd1 vccd1 vccd1 _09380_ sky130_fd_sc_hd__nand3_1
X_19526_ _03000_ _03001_ _03002_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19457_ rbzero.debug_overlay.vplaneY\[0\] rbzero.debug_overlay.vplaneY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__and2_1
X_16669_ _09309_ _09310_ _09266_ vssd1 vssd1 vccd1 vccd1 _09312_ sky130_fd_sc_hd__a21o_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18408_ _01965_ _01929_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__or2b_1
XFILLER_34_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19388_ _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__nand2_1
XFILLER_195_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18339_ _02036_ _02037_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__nand2_1
XFILLER_147_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21350_ net271 _01119_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21281_ clknet_leaf_37_i_clk _01050_ vssd1 vssd1 vccd1 vccd1 rbzero.hsync sky130_fd_sc_hd__dfxtp_1
XFILLER_190_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20094_ clknet_1_0__leaf__03044_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__buf_1
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_54_i_clk clknet_3_7_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19631__83 clknet_1_1__leaf__03043_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__inv_2
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20996_ clknet_leaf_10_i_clk _00765_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1067 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10680_ rbzero.tex_g1\[17\] rbzero.tex_g1\[18\] _03680_ vssd1 vssd1 vccd1 vccd1 _03681_
+ sky130_fd_sc_hd__mux2_1
XFILLER_111_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21617_ clknet_leaf_27_i_clk _01386_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12350_ _04813_ _04811_ _04006_ _03475_ _05083_ _05082_ vssd1 vssd1 vccd1 vccd1 _05118_
+ sky130_fd_sc_hd__mux4_1
X_21548_ net469 _01317_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11301_ _04077_ _04080_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__nor2_1
X_12281_ _04021_ _05047_ _05049_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__and3_1
XFILLER_181_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21479_ net400 _01248_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_135_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14020_ _06755_ _06756_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__nor2_1
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11232_ _04016_ _03997_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__or2_2
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11163_ _03946_ _03949_ _03950_ _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__or4_1
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11094_ _03897_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__clkbuf_1
X_15971_ _08584_ _08614_ _08615_ vssd1 vssd1 vccd1 vccd1 _08616_ sky130_fd_sc_hd__a21oi_4
XFILLER_150_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17710_ _10122_ _10146_ _10274_ vssd1 vssd1 vccd1 vccd1 _10275_ sky130_fd_sc_hd__a21o_1
X_14922_ rbzero.wall_tracer.trackDistY\[-1\] rbzero.wall_tracer.trackDistX\[-1\] _07616_
+ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__mux2_1
X_18690_ _02383_ _02385_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__xnor2_2
XFILLER_121_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ _09526_ _09029_ _09165_ _09245_ vssd1 vssd1 vccd1 vccd1 _10206_ sky130_fd_sc_hd__o22a_1
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ rbzero.wall_tracer.stepDistY\[6\] _07571_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07572_ sky130_fd_sc_hd__mux2_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ _06534_ _06538_ _06539_ _06540_ _06518_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__a311o_1
XFILLER_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17572_ rbzero.wall_tracer.stepDistX\[10\] vssd1 vssd1 vccd1 vccd1 _10138_ sky130_fd_sc_hd__inv_2
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14784_ _07498_ _07489_ _05952_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__mux2_1
XFILLER_147_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11996_ _04232_ _04758_ _04762_ _04770_ _04244_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__o311a_1
XFILLER_95_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19311_ _02811_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_204_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16523_ _09033_ _09035_ _09032_ vssd1 vssd1 vccd1 vccd1 _09167_ sky130_fd_sc_hd__a21bo_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13735_ _06382_ _06153_ _06469_ _06470_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__a22o_1
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10947_ rbzero.tex_b1\[18\] rbzero.tex_b1\[19\] _03817_ vssd1 vssd1 vccd1 vccd1 _03821_
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19242_ _02561_ _02772_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__or2_1
XFILLER_177_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16454_ _09095_ _09097_ vssd1 vssd1 vccd1 vccd1 _09098_ sky130_fd_sc_hd__and2_1
X_13666_ _06356_ _06401_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ rbzero.tex_b1\[51\] rbzero.tex_b1\[52\] _03784_ vssd1 vssd1 vccd1 vccd1 _03785_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15405_ rbzero.wall_tracer.side rbzero.wall_tracer.rayAddendX\[-2\] vssd1 vssd1 vccd1
+ vccd1 _08050_ sky130_fd_sc_hd__nand2_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19173_ _05190_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__buf_4
X_12617_ _05324_ _05325_ _05326_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__a21bo_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _09029_ _08162_ vssd1 vssd1 vccd1 vccd1 _09030_ sky130_fd_sc_hd__nor2_2
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13597_ _06279_ _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__and2_1
X_18124_ _09391_ _09703_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__and2_1
XFILLER_118_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15336_ _07980_ vssd1 vssd1 vccd1 vccd1 _07981_ sky130_fd_sc_hd__clkbuf_4
X_12548_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__nor2_1
XFILLER_172_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18055_ _08895_ _01524_ _10266_ _08767_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__o22ai_1
XFILLER_32_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15267_ _05206_ _07902_ _07910_ _07911_ vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__a22o_4
XANTENNA_2 _05190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _05233_ _05216_ _05213_ _05230_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__or4_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17006_ _09640_ _09645_ vssd1 vssd1 vccd1 vccd1 _09646_ sky130_fd_sc_hd__xnor2_1
X_14218_ _06892_ _06954_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__xnor2_1
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15198_ _07849_ _07850_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__nand2_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14149_ _06860_ _06874_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__xnor2_1
XFILLER_99_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20210__233 clknet_1_1__leaf__03303_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__inv_2
XFILLER_140_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18957_ _02608_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17908_ _01609_ _01610_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__and2_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18888_ rbzero.spi_registers.sclk_buffer\[2\] rbzero.spi_registers.sclk_buffer\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__nor2b_2
XFILLER_6_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17839_ _01454_ _01542_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__xnor2_1
XFILLER_82_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20850_ clknet_leaf_44_i_clk _00619_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19509_ _03913_ _02986_ _02987_ _07855_ rbzero.wall_tracer.rayAddendY\[7\] vssd1
+ vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__a32o_1
XFILLER_63_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20781_ clknet_leaf_72_i_clk _00550_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21402_ net323 _01171_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21333_ net254 _01102_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21264_ clknet_leaf_97_i_clk _01033_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-2\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_2_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21195_ clknet_leaf_92_i_clk _00964_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20185__210 clknet_1_1__leaf__03301_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__inv_2
XFILLER_131_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _04244_ _04618_ _04626_ _04116_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a31o_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _03744_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _04557_ _04558_ _04218_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__mux2_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20979_ clknet_leaf_8_i_clk _00748_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_202_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13520_ _06214_ _06217_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__and2b_1
X_10732_ rbzero.tex_g0\[57\] rbzero.tex_g0\[56\] _03706_ vssd1 vssd1 vccd1 vccd1 _03708_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13451_ _06172_ _06187_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__xnor2_1
X_10663_ rbzero.tex_g1\[25\] rbzero.tex_g1\[26\] _03669_ vssd1 vssd1 vccd1 vccd1 _03672_
+ sky130_fd_sc_hd__mux2_1
XFILLER_90_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12402_ _04813_ _04811_ _05143_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__mux2_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16170_ _08813_ _08814_ vssd1 vssd1 vccd1 vccd1 _08815_ sky130_fd_sc_hd__or2_1
X_10594_ _03482_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__clkbuf_4
XFILLER_142_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13382_ _05923_ _06116_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__nand2_1
XFILLER_182_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15121_ _07754_ _07763_ _07764_ _07749_ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__o2bb2ai_1
X_12333_ _05100_ net28 vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__nand2_1
XFILLER_5_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15052_ _07712_ _07714_ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__xnor2_1
X_12264_ net22 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__inv_2
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14003_ _06739_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__clkbuf_4
X_11215_ rbzero.wall_tracer.state\[11\] vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__inv_2
X_12195_ _04962_ _04963_ _04964_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__and3_1
X_19860_ rbzero.debug_overlay.playerX\[1\] _03167_ vssd1 vssd1 vccd1 vccd1 _03172_
+ sky130_fd_sc_hd__and2_1
XFILLER_107_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput61 net61 vssd1 vssd1 vccd1 vccd1 o_rgb[14] sky130_fd_sc_hd__buf_2
X_18811_ _05254_ _08186_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__nor2_1
X_11146_ rbzero.map_rom.i_row\[4\] vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__clkinv_2
XFILLER_150_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19791_ _03124_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18742_ _02428_ _02429_ _02430_ _05531_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a31o_1
X_11077_ rbzero.tex_b0\[21\] rbzero.tex_b0\[20\] _03887_ vssd1 vssd1 vccd1 vccd1 _03889_
+ sky130_fd_sc_hd__mux2_1
X_15954_ _08590_ _08597_ vssd1 vssd1 vccd1 vccd1 _08599_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__03291_ clknet_0__03291_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03291_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_110_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14905_ _07591_ _07610_ _07611_ _04039_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__o211a_1
X_18673_ _01737_ _01524_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__or2_1
XFILLER_48_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15885_ _08526_ _08528_ _08529_ vssd1 vssd1 vccd1 vccd1 _08530_ sky130_fd_sc_hd__a21oi_2
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17624_ _10064_ _10067_ _10188_ vssd1 vssd1 vccd1 vccd1 _10189_ sky130_fd_sc_hd__a21o_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14836_ _07559_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__clkbuf_4
XFILLER_184_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19610__64 clknet_1_1__leaf__03041_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__inv_2
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17555_ _10119_ _10120_ vssd1 vssd1 vccd1 vccd1 _10121_ sky130_fd_sc_hd__or2b_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14767_ _05814_ _07496_ _07500_ _07486_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__a211oi_1
X_11979_ _04242_ _04745_ _04753_ _04207_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__o211a_1
X_16506_ _08991_ _08993_ vssd1 vssd1 vccd1 vccd1 _09150_ sky130_fd_sc_hd__or2b_1
XFILLER_205_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_204_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13718_ _06439_ _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__xor2_1
XFILLER_108_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17486_ _09971_ _09957_ vssd1 vssd1 vccd1 vccd1 _10052_ sky130_fd_sc_hd__or2b_1
XFILLER_177_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14698_ _07106_ _07419_ _07420_ _07423_ _05892_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__a311o_1
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19225_ rbzero.spi_registers.got_new_vshift _02711_ vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__nand2_2
X_16437_ _09081_ vssd1 vssd1 vccd1 vccd1 _09082_ sky130_fd_sc_hd__buf_4
XFILLER_108_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ _06339_ _06383_ _06384_ _06385_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19156_ rbzero.otherx\[4\] _02710_ _02718_ _02714_ vssd1 vssd1 vccd1 vccd1 _00733_
+ sky130_fd_sc_hd__o211a_1
X_16368_ _09011_ _09012_ vssd1 vssd1 vccd1 vccd1 _09013_ sky130_fd_sc_hd__xnor2_1
XFILLER_121_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18107_ _01701_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__inv_2
XFILLER_8_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15319_ _04013_ _07962_ _07963_ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__a21oi_4
XFILLER_184_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19087_ rbzero.spi_registers.spi_counter\[3\] rbzero.spi_registers.spi_counter\[2\]
+ _02567_ _02558_ _02557_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__o311a_1
X_16299_ _08764_ _08807_ _08811_ _08940_ _08943_ vssd1 vssd1 vccd1 vccd1 _08944_ sky130_fd_sc_hd__a32oi_4
X_18038_ _01739_ _10238_ _09552_ _01737_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__o22ai_1
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20000_ rbzero.pov.ready_buffer\[4\] _03246_ _03248_ rbzero.debug_overlay.vplaneY\[-5\]
+ _02741_ vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__a221o_1
XFILLER_113_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19989_ rbzero.pov.ready_buffer\[15\] _03246_ _03248_ rbzero.debug_overlay.vplaneX\[-5\]
+ _03251_ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__a221o_1
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ clknet_leaf_87_i_clk _00671_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20833_ clknet_leaf_54_i_clk _00602_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20764_ clknet_leaf_45_i_clk _00533_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20695_ clknet_leaf_58_i_clk _00479_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20217__239 clknet_1_0__leaf__03304_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__inv_2
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21316_ net237 _01085_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21247_ clknet_leaf_91_i_clk _01016_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_85_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11000_ _03848_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21178_ clknet_leaf_5_i_clk _00947_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12951_ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__inv_2
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ rbzero.tex_b0\[3\] _04135_ _04136_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__and3_1
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15670_ _07959_ _07941_ vssd1 vssd1 vccd1 vccd1 _08315_ sky130_fd_sc_hd__nor2_1
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12882_ _05610_ _05612_ _05615_ _05601_ _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__a2111o_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _07316_ _07317_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__xnor2_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _04242_ _04601_ _04609_ _04207_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__o211a_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17340_ _09486_ _09495_ vssd1 vssd1 vccd1 vccd1 _09907_ sky130_fd_sc_hd__and2b_1
XFILLER_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _07058_ _06999_ _07000_ _07057_ _07055_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__o32ai_2
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _04540_ _04541_ _04126_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__mux2_1
XFILLER_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13503_ _06159_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__clkbuf_4
XFILLER_41_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ rbzero.tex_g1\[0\] rbzero.tex_g1\[1\] _03691_ vssd1 vssd1 vccd1 vccd1 _03699_
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _09845_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14483_ _07168_ _07219_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__nand2_1
X_11695_ rbzero.debug_overlay.vplaneY\[-7\] _04455_ _04465_ rbzero.debug_overlay.vplaneY\[-1\]
+ _04040_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__a221o_1
X_19010_ rbzero.pov.spi_buffer\[37\] rbzero.pov.ready_buffer\[37\] _02627_ vssd1 vssd1
+ vccd1 vccd1 _02636_ sky130_fd_sc_hd__mux2_1
XFILLER_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16222_ _08865_ _08866_ vssd1 vssd1 vccd1 vccd1 _08867_ sky130_fd_sc_hd__and2_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13434_ _06004_ _06005_ _06019_ _06020_ _06001_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__a32o_1
X_10646_ rbzero.tex_g1\[33\] rbzero.tex_g1\[34\] _03658_ vssd1 vssd1 vccd1 vccd1 _03663_
+ sky130_fd_sc_hd__mux2_1
XFILLER_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ _08779_ _08797_ vssd1 vssd1 vccd1 vccd1 _08798_ sky130_fd_sc_hd__nand2_1
X_13365_ _06100_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__or2_1
XFILLER_182_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10577_ _03626_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__clkbuf_1
X_20157__186 clknet_1_1__leaf__03297_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__inv_2
X_15104_ _04462_ rbzero.debug_overlay.vplaneX\[-7\] vssd1 vssd1 vccd1 vccd1 _07763_
+ sky130_fd_sc_hd__xnor2_1
X_12316_ _05082_ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__nor2_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16084_ _07912_ _08125_ vssd1 vssd1 vccd1 vccd1 _08729_ sky130_fd_sc_hd__or2_1
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ _05939_ _05975_ _05962_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__or3b_1
XFILLER_108_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15035_ _07680_ _07693_ _07681_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__o21ai_1
X_19912_ rbzero.pov.ready_buffer\[51\] _02823_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__nand2_1
X_12247_ _04996_ _05013_ _05016_ net16 vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__o22a_1
XFILLER_123_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19843_ _03139_ _03158_ _03159_ _03157_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__o211a_1
X_12178_ _04883_ _04884_ gpout0.vpos\[6\] _04887_ _04910_ net10 vssd1 vssd1 vccd1
+ vccd1 _04949_ sky130_fd_sc_hd__mux4_1
X_11129_ rbzero.wall_tracer.visualWallDist\[10\] rbzero.wall_tracer.visualWallDist\[9\]
+ _03916_ _03917_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__or4_1
X_19774_ rbzero.pov.spi_buffer\[60\] rbzero.pov.spi_buffer\[61\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03116_ sky130_fd_sc_hd__mux2_1
X_16986_ _09624_ _09625_ vssd1 vssd1 vccd1 vccd1 _09626_ sky130_fd_sc_hd__and2_1
XFILLER_77_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18725_ _02414_ _02415_ _02416_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__and3_1
X_15937_ _08578_ _08580_ _08581_ vssd1 vssd1 vccd1 vccd1 _08582_ sky130_fd_sc_hd__o21ai_2
XFILLER_3_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18656_ _02247_ _02236_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__and2b_1
X_15868_ _08456_ _08457_ vssd1 vssd1 vccd1 vccd1 _08513_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20322__334 clknet_1_1__leaf__03314_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__inv_2
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14819_ rbzero.wall_tracer.stepDistY\[-3\] _07545_ _07546_ vssd1 vssd1 vccd1 vccd1
+ _07547_ sky130_fd_sc_hd__mux2_1
X_17607_ _10172_ vssd1 vssd1 vccd1 vccd1 _10173_ sky130_fd_sc_hd__inv_2
X_18587_ _02282_ _02283_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__nor2_1
XFILLER_52_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15799_ _08379_ _08443_ vssd1 vssd1 vccd1 vccd1 _08444_ sky130_fd_sc_hd__xor2_2
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17538_ _09670_ _09964_ vssd1 vssd1 vccd1 vccd1 _10104_ sky130_fd_sc_hd__nand2_1
XFILLER_33_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17469_ _09817_ vssd1 vssd1 vccd1 vccd1 _10036_ sky130_fd_sc_hd__buf_2
XFILLER_178_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19208_ rbzero.spi_registers.new_floor\[0\] rbzero.color_floor\[0\] _02751_ vssd1
+ vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__mux2_1
XFILLER_34_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20480_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__inv_2
XFILLER_177_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19139_ _04037_ _02705_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__nand2_1
XFILLER_157_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21101_ net191 _00870_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[41\] sky130_fd_sc_hd__dfxtp_1
XFILLER_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21032_ clknet_leaf_13_i_clk _00801_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20297__311 clknet_1_0__leaf__03312_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__inv_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20816_ clknet_leaf_58_i_clk _00585_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20747_ clknet_leaf_39_i_clk _00516_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_204_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10500_ rbzero.tex_r0\[39\] rbzero.tex_r0\[38\] _03580_ vssd1 vssd1 vccd1 vccd1 _03586_
+ sky130_fd_sc_hd__mux2_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11480_ _04219_ _04259_ _04254_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__o21a_1
XFILLER_168_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20678_ clknet_leaf_49_i_clk _00462_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[7\]
+ sky130_fd_sc_hd__dfxtp_4
Xclkbuf_1_0__f__03294_ clknet_0__03294_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03294_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_195_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10431_ _03547_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13150_ _05883_ _05886_ _05798_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__o21a_1
X_10362_ _03511_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_136_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12101_ _04317_ _04853_ _04838_ _03473_ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__a221o_1
XFILLER_191_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13081_ _05690_ _05796_ _05817_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__o21a_1
XFILLER_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12032_ _04805_ _04806_ _04206_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__mux2_1
XFILLER_151_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16840_ rbzero.wall_tracer.visualWallDist\[10\] _04015_ vssd1 vssd1 vccd1 vccd1 _09481_
+ sky130_fd_sc_hd__nand2_2
XFILLER_120_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16771_ _09411_ _09412_ vssd1 vssd1 vccd1 vccd1 _09413_ sky130_fd_sc_hd__xor2_2
XFILLER_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13983_ _06674_ _06679_ _06673_ _06683_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__a22oi_2
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18510_ _02078_ _02081_ _02207_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__a21o_1
X_15722_ _08350_ _08351_ _08366_ vssd1 vssd1 vccd1 vccd1 _08367_ sky130_fd_sc_hd__a21o_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12934_ _05563_ _05653_ _05669_ _05650_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__a211o_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _02968_ _02969_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__xor2_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18441_ _02028_ _01645_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__and2b_1
X_15653_ _08262_ _08278_ vssd1 vssd1 vccd1 vccd1 _08298_ sky130_fd_sc_hd__xnor2_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12865_ rbzero.wall_tracer.visualWallDist\[5\] _04031_ vssd1 vssd1 vccd1 vccd1 _05602_
+ sky130_fd_sc_hd__nor2_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20163__190 clknet_1_0__leaf__03299_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__inv_2
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14604_ _07206_ _07339_ _07338_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__or3_1
XFILLER_61_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _01498_ _09162_ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__nor2_1
X_11816_ _04591_ _04593_ _04324_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__o21ba_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15584_ _08216_ _08228_ vssd1 vssd1 vccd1 vccd1 _08229_ sky130_fd_sc_hd__xnor2_4
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _05533_ _05537_ _05538_ _05284_ rbzero.wall_tracer.mapY\[6\] vssd1 vssd1
+ vccd1 vccd1 _00413_ sky130_fd_sc_hd__a32o_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _09880_ _09882_ _09881_ vssd1 vssd1 vccd1 vccd1 _09892_ sky130_fd_sc_hd__a21boi_1
XFILLER_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _07252_ _07267_ _07271_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__o21a_1
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ rbzero.tex_g0\[13\] rbzero.tex_g0\[12\] _04271_ vssd1 vssd1 vccd1 vccd1 _04525_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17254_ rbzero.wall_tracer.trackDistX\[-9\] rbzero.wall_tracer.stepDistX\[-9\] vssd1
+ vssd1 vccd1 vccd1 _09830_ sky130_fd_sc_hd__or2_1
XFILLER_187_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14466_ _07132_ _07201_ _07202_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__o21ai_1
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ rbzero.debug_overlay.vplaneX\[-5\] _04454_ _04455_ rbzero.debug_overlay.vplaneX\[-7\]
+ _04456_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__a221o_1
X_16205_ _08845_ _08847_ _08849_ vssd1 vssd1 vccd1 vccd1 _08850_ sky130_fd_sc_hd__a21o_1
X_13417_ _05752_ _06153_ _05976_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__and3_1
X_10629_ rbzero.tex_g1\[41\] rbzero.tex_g1\[42\] _03647_ vssd1 vssd1 vccd1 vccd1 _03654_
+ sky130_fd_sc_hd__mux2_1
X_17185_ rbzero.wall_tracer.wall\[0\] rbzero.row_render.wall\[0\] _07830_ vssd1 vssd1
+ vccd1 vccd1 _09772_ sky130_fd_sc_hd__mux2_1
X_14397_ _07114_ _07127_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__nand2_1
XFILLER_183_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16136_ _08743_ _08750_ vssd1 vssd1 vccd1 vccd1 _08781_ sky130_fd_sc_hd__or2_1
X_13348_ _06041_ _06084_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__nor2_1
XFILLER_115_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16067_ _08698_ _08711_ vssd1 vssd1 vccd1 vccd1 _08712_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13279_ _06011_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15018_ rbzero.debug_overlay.vplaneX\[-6\] rbzero.wall_tracer.rayAddendX\[-6\] vssd1
+ vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__or2_1
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19826_ rbzero.pov.ready_buffer\[60\] _07985_ _03146_ vssd1 vssd1 vccd1 vccd1 _03147_
+ sky130_fd_sc_hd__mux2_1
XFILLER_190_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19757_ rbzero.pov.spi_buffer\[52\] rbzero.pov.spi_buffer\[53\] _03103_ vssd1 vssd1
+ vccd1 vccd1 _03107_ sky130_fd_sc_hd__mux2_1
XFILLER_96_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16969_ _09485_ _09486_ _09497_ _09608_ vssd1 vssd1 vccd1 vccd1 _09609_ sky130_fd_sc_hd__a31o_1
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18708_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__nand2_1
X_19688_ rbzero.pov.spi_buffer\[19\] rbzero.pov.spi_buffer\[20\] _03070_ vssd1 vssd1
+ vccd1 vccd1 _03071_ sky130_fd_sc_hd__mux2_1
XFILLER_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18639_ _02333_ _02334_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__xnor2_1
XFILLER_25_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21650_ clknet_leaf_43_i_clk _01419_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texVinit\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20601_ gpout2.clk_div\[0\] gpout2.clk_div\[1\] vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__nand2_1
XFILLER_36_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21581_ net502 _01350_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20532_ rbzero.traced_texa\[8\] rbzero.texV\[8\] vssd1 vssd1 vccd1 vccd1 _03424_
+ sky130_fd_sc_hd__nor2_1
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20463_ _03272_ _03365_ _03366_ _03327_ rbzero.texV\[-4\] vssd1 vssd1 vccd1 vccd1
+ _01392_ sky130_fd_sc_hd__a32o_1
XFILLER_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21015_ clknet_leaf_8_i_clk _00784_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_101_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10980_ rbzero.tex_b1\[2\] rbzero.tex_b1\[3\] _03828_ vssd1 vssd1 vccd1 vccd1 _03838_
+ sky130_fd_sc_hd__mux2_1
XFILLER_83_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12650_ _05398_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11601_ rbzero.tex_r1\[56\] _04273_ _04379_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__a21o_1
XFILLER_90_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _05333_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__or2_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14320_ _07013_ _07014_ _07056_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__o21a_1
XFILLER_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11532_ rbzero.color_sky\[0\] rbzero.color_floor\[0\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04312_ sky130_fd_sc_hd__mux2_2
XFILLER_184_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ _06986_ _06987_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__xnor2_1
XFILLER_183_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11463_ _04230_ _04236_ _04240_ _04242_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__a211o_1
XFILLER_139_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13202_ _05938_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__buf_4
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10414_ rbzero.tex_r1\[13\] rbzero.tex_r1\[14\] _03538_ vssd1 vssd1 vccd1 vccd1 _03539_
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14182_ _06709_ _06918_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__nand2_1
XFILLER_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11394_ gpout0.hpos\[7\] _04159_ _04157_ gpout0.hpos\[8\] _04173_ vssd1 vssd1 vccd1
+ vccd1 _04174_ sky130_fd_sc_hd__o221a_1
XFILLER_48_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20351__360 clknet_1_0__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__inv_2
XFILLER_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ _05820_ _05866_ _05869_ _05813_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__o211a_1
XFILLER_174_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10345_ _03502_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__clkbuf_1
X_18990_ _02625_ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17941_ _01641_ _01642_ _01634_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__a21o_1
XFILLER_124_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _05796_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__clkbuf_4
XFILLER_79_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12015_ _04788_ _04789_ _04304_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__mux2_1
XFILLER_78_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17872_ _01494_ _01512_ _01574_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__a21oi_1
X_20269__287 clknet_1_1__leaf__03308_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__inv_2
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16823_ _09463_ _09464_ vssd1 vssd1 vccd1 vccd1 _09465_ sky130_fd_sc_hd__nor2_1
XFILLER_94_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19542_ _07677_ _03016_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__nor2_1
X_16754_ _08111_ _08264_ vssd1 vssd1 vccd1 vccd1 _09396_ sky130_fd_sc_hd__and2b_1
X_13966_ _06685_ _06695_ _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15705_ _08320_ _08322_ vssd1 vssd1 vccd1 vccd1 _08350_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1__f__03042_ clknet_0__03042_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03042_
+ sky130_fd_sc_hd__clkbuf_16
X_12917_ _05563_ _05653_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__nand2_1
X_16685_ _09208_ _09327_ vssd1 vssd1 vccd1 vccd1 _09328_ sky130_fd_sc_hd__nand2_1
X_19473_ _02951_ _02952_ _02950_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a21o_1
X_13897_ _06632_ _06633_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__and2_1
XFILLER_185_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18424_ _02009_ _01917_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__or2b_1
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15636_ _08249_ _08280_ vssd1 vssd1 vccd1 vccd1 _08281_ sky130_fd_sc_hd__xor2_4
X_12848_ rbzero.wall_tracer.visualWallDist\[-6\] rbzero.wall_tracer.rcp_sel\[2\] vssd1
+ vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or2_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18355_ _02038_ _02053_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__xnor2_1
X_15567_ _07894_ _05331_ _08211_ _07970_ vssd1 vssd1 vccd1 vccd1 _08212_ sky130_fd_sc_hd__o211a_1
XFILLER_148_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ rbzero.map_rom.i_col\[4\] _05523_ _05414_ vssd1 vssd1 vccd1 vccd1 _05524_
+ sky130_fd_sc_hd__mux2_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14518_ _07230_ _07229_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__and2b_1
X_17306_ _09807_ _09331_ vssd1 vssd1 vccd1 vccd1 _09877_ sky130_fd_sc_hd__or2_1
XFILLER_159_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18286_ _01860_ _01620_ _01984_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__o21ai_1
X_15498_ _08138_ _08142_ vssd1 vssd1 vccd1 vccd1 _08143_ sky130_fd_sc_hd__xor2_1
XFILLER_70_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14449_ _07114_ _07185_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__nor2_1
X_17237_ rbzero.wall_tracer.trackDistX\[-12\] rbzero.wall_tracer.stepDistX\[-12\]
+ _09813_ _09814_ vssd1 vssd1 vccd1 vccd1 _09815_ sky130_fd_sc_hd__and4_1
XFILLER_128_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17168_ _07679_ vssd1 vssd1 vccd1 vccd1 _09769_ sky130_fd_sc_hd__clkbuf_4
XFILLER_190_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16119_ _08719_ _08763_ vssd1 vssd1 vccd1 vccd1 _08764_ sky130_fd_sc_hd__xor2_2
XFILLER_192_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17099_ _09737_ _09738_ vssd1 vssd1 vccd1 vccd1 _09739_ sky130_fd_sc_hd__xnor2_4
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19809_ _03133_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03309_ clknet_0__03309_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03309_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_opt_8_0_i_clk clknet_3_3_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_8_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_197_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21633_ clknet_leaf_32_i_clk _01402_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21564_ net485 _01333_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20515_ rbzero.texV\[4\] _03327_ _03332_ _03410_ vssd1 vssd1 vccd1 vccd1 _01400_
+ sky130_fd_sc_hd__a22o_1
X_21495_ net416 _01264_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_181_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20446_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1 _03352_
+ sky130_fd_sc_hd__nand2_1
XFILLER_107_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13820_ _06279_ _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__xnor2_2
XFILLER_75_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13751_ _06486_ _06487_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__nand2_1
X_10963_ _03829_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_204_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12702_ _05446_ _05447_ _05449_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__o21a_1
XFILLER_203_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16470_ _07959_ vssd1 vssd1 vccd1 vccd1 _09114_ sky130_fd_sc_hd__clkbuf_4
X_13682_ _06393_ _06418_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__xnor2_1
XFILLER_188_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10894_ rbzero.tex_b1\[43\] rbzero.tex_b1\[44\] _03784_ vssd1 vssd1 vccd1 vccd1 _03793_
+ sky130_fd_sc_hd__mux2_1
XFILLER_188_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15421_ _08027_ _08065_ vssd1 vssd1 vccd1 vccd1 _08066_ sky130_fd_sc_hd__nand2_1
X_12633_ rbzero.debug_overlay.playerY\[2\] _05385_ _05204_ vssd1 vssd1 vccd1 vccd1
+ _05386_ sky130_fd_sc_hd__mux2_1
XFILLER_19_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18140_ _01498_ _01475_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__nor2_1
XFILLER_169_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15352_ _07977_ _07981_ _07989_ _07996_ vssd1 vssd1 vccd1 vccd1 _07997_ sky130_fd_sc_hd__o22ai_1
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12564_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__inv_2
XFILLER_180_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14303_ _07035_ _07038_ _07039_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__nor3b_2
XFILLER_106_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18071_ _01770_ _01771_ _01772_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__nand3_1
X_11515_ rbzero.tex_r0\[21\] rbzero.tex_r0\[20\] _04291_ vssd1 vssd1 vccd1 vccd1 _04295_
+ sky130_fd_sc_hd__mux2_1
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15283_ _07904_ rbzero.wall_tracer.stepDistY\[-4\] _05195_ vssd1 vssd1 vccd1 vccd1
+ _07928_ sky130_fd_sc_hd__a21o_1
X_12495_ rbzero.wall_tracer.trackDistY\[-5\] _05236_ rbzero.wall_tracer.trackDistY\[-6\]
+ _05237_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__o221a_1
XFILLER_106_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17022_ _08204_ _09103_ _08493_ _08383_ vssd1 vssd1 vccd1 vccd1 _09662_ sky130_fd_sc_hd__o22ai_1
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20275__291 clknet_1_1__leaf__03310_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__inv_2
XFILLER_144_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14234_ _06805_ _06678_ _06937_ vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__o21bai_1
X_11446_ _04225_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__clkbuf_4
XFILLER_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14165_ _06680_ _06690_ _06672_ _06675_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__o22a_1
X_11377_ _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__and2_1
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13116_ _05794_ _05828_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__or2_2
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10328_ _03493_ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__clkbuf_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _06826_ _06831_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__nor2_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ rbzero.pov.spi_buffer\[19\] rbzero.pov.ready_buffer\[19\] _02616_ vssd1 vssd1
+ vccd1 vccd1 _02617_ sky130_fd_sc_hd__mux2_1
XFILLER_112_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _10244_ _01503_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__nand2_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _05719_ _05721_ _05705_ _05783_ _05710_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__o32a_1
XFILLER_61_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17855_ _09889_ _01558_ _09781_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16806_ _09382_ _09447_ vssd1 vssd1 vccd1 vccd1 _09448_ sky130_fd_sc_hd__xnor2_1
X_17786_ _01471_ _01489_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__xor2_1
X_14998_ _07669_ vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_47_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19525_ _02906_ rbzero.wall_tracer.rayAddendY\[9\] vssd1 vssd1 vccd1 vccd1 _03002_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_75_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16737_ _09263_ _09349_ _09378_ vssd1 vssd1 vccd1 vccd1 _09379_ sky130_fd_sc_hd__a21o_1
XFILLER_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13949_ _06665_ _06670_ _06684_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__nand3_1
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19456_ rbzero.debug_overlay.vplaneY\[0\] rbzero.debug_overlay.vplaneY\[-4\] vssd1
+ vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__nor2_1
XFILLER_62_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16668_ _09266_ _09309_ _09310_ vssd1 vssd1 vccd1 vccd1 _09311_ sky130_fd_sc_hd__nand3_1
XFILLER_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18407_ _01964_ _01932_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__or2b_1
X_15619_ _08199_ _08201_ _08203_ vssd1 vssd1 vccd1 vccd1 _08264_ sky130_fd_sc_hd__a21bo_2
X_19387_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__nand2_1
X_16599_ _09124_ _09116_ vssd1 vssd1 vccd1 vccd1 _09242_ sky130_fd_sc_hd__or2b_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18338_ _01971_ _01968_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__or2b_1
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18269_ _10110_ _01524_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__nor2_1
XFILLER_190_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21280_ clknet_leaf_36_i_clk _01049_ vssd1 vssd1 vccd1 vccd1 rbzero.vga_sync.vsync
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_190_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20995_ clknet_leaf_1_i_clk _00764_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.spi_done
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21616_ clknet_leaf_27_i_clk _01385_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_187_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21547_ net468 _01316_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ rbzero.texV\[3\] _04078_ _04079_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__a21boi_1
X_12280_ net21 net20 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__and2_1
X_21478_ net399 _01247_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11231_ rbzero.wall_tracer.state\[1\] vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__clkinv_4
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20429_ rbzero.traced_texa\[-9\] rbzero.texV\[-9\] vssd1 vssd1 vccd1 vccd1 _03338_
+ sky130_fd_sc_hd__or2_1
XFILLER_150_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__03045_ clknet_0__03045_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03045_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11162_ rbzero.wall_tracer.mapX\[11\] rbzero.wall_tracer.mapX\[10\] rbzero.wall_tracer.mapY\[7\]
+ rbzero.wall_tracer.mapY\[6\] vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__or4_1
XFILLER_107_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15970_ _08585_ _08613_ vssd1 vssd1 vccd1 vccd1 _08615_ sky130_fd_sc_hd__nor2_1
XFILLER_1_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11093_ rbzero.tex_b0\[13\] rbzero.tex_b0\[12\] _03887_ vssd1 vssd1 vccd1 vccd1 _03897_
+ sky130_fd_sc_hd__mux2_1
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14921_ _07621_ _07622_ _07623_ _07620_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__o211a_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ _08705_ _09029_ _09165_ vssd1 vssd1 vccd1 vccd1 _10205_ sky130_fd_sc_hd__or3_1
X_14852_ _07394_ _07433_ _07418_ _07468_ _07570_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__a311o_4
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13803_ _06503_ _06516_ _06517_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__a21oi_1
X_17571_ _09117_ _09977_ vssd1 vssd1 vccd1 vccd1 _10137_ sky130_fd_sc_hd__nor2_1
X_14783_ _00004_ _07514_ _07515_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a21oi_1
XFILLER_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11995_ _04306_ _04765_ _04769_ _04241_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__a211o_1
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19310_ rbzero.spi_registers.new_other\[10\] rbzero.spi_registers.spi_buffer\[10\]
+ _02800_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__mux2_1
X_16522_ _09029_ _08160_ _09165_ _08162_ vssd1 vssd1 vccd1 vccd1 _09166_ sky130_fd_sc_hd__o22a_1
XFILLER_147_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13734_ _06382_ _06153_ _06469_ _06470_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__nand4_1
XFILLER_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10946_ _03820_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_205_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19241_ rbzero.spi_registers.spi_done _03480_ _02560_ vssd1 vssd1 vccd1 vccd1 _02772_
+ sky130_fd_sc_hd__nand3_1
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16453_ _09096_ _08356_ _09094_ vssd1 vssd1 vccd1 vccd1 _09097_ sky130_fd_sc_hd__o21ai_1
X_13665_ _06041_ _06016_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__or2_1
XFILLER_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10877_ _03646_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ _05342_ _05345_ _05365_ _05369_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or4b_2
X_15404_ rbzero.wall_tracer.rayAddendY\[-2\] vssd1 vssd1 vccd1 vccd1 _08049_ sky130_fd_sc_hd__inv_2
X_16384_ _09028_ vssd1 vssd1 vccd1 vccd1 _09029_ sky130_fd_sc_hd__clkbuf_4
X_19172_ rbzero.spi_registers.got_new_vinf _02711_ rbzero.row_render.vinf vssd1 vssd1
+ vccd1 vccd1 _02729_ sky130_fd_sc_hd__a21o_1
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13596_ _06331_ _06332_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__and2b_1
XFILLER_197_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18123_ _01822_ _01823_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__or2_1
XFILLER_157_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15335_ rbzero.debug_overlay.playerX\[-9\] _05206_ _07979_ vssd1 vssd1 vccd1 vccd1
+ _07980_ sky130_fd_sc_hd__a21oi_4
X_12547_ rbzero.debug_overlay.facingY\[-5\] rbzero.wall_tracer.rayAddendY\[3\] vssd1
+ vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__and2_1
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18054_ _10131_ _10132_ _01525_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__a21o_2
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15266_ rbzero.wall_tracer.visualWallDist\[-6\] _04013_ _05195_ vssd1 vssd1 vccd1
+ vccd1 _07911_ sky130_fd_sc_hd__a21oi_1
X_12478_ _05219_ _05221_ _05223_ _05225_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__or4_1
XFILLER_32_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_3 _05204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17005_ _09641_ _09644_ vssd1 vssd1 vccd1 vccd1 _09645_ sky130_fd_sc_hd__xnor2_1
X_14217_ _06900_ _06899_ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__and2b_1
XFILLER_126_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11429_ _04208_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__buf_6
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15197_ _07730_ _07833_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__nand2_1
XFILLER_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14148_ _06858_ _06876_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__xnor2_1
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14079_ _06799_ _06814_ _06815_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__a21bo_1
X_18956_ rbzero.pov.spi_buffer\[11\] rbzero.pov.ready_buffer\[11\] _02605_ vssd1 vssd1
+ vccd1 vccd1 _02608_ sky130_fd_sc_hd__mux2_1
XFILLER_100_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17907_ _01573_ _01608_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__or2_1
XFILLER_117_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18887_ rbzero.spi_registers.ss_buffer\[1\] _03555_ vssd1 vssd1 vccd1 vccd1 _02557_
+ sky130_fd_sc_hd__nor2_2
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17838_ _01539_ _01541_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__xor2_1
XFILLER_187_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17769_ _10240_ _10242_ _10237_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__a21bo_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19508_ _02984_ _02985_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__or2_1
XFILLER_74_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20780_ clknet_leaf_72_i_clk _00549_ vssd1 vssd1 vccd1 vccd1 rbzero.traced_texa\[-8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19439_ rbzero.debug_overlay.vplaneY\[10\] rbzero.wall_tracer.rayAddendY\[2\] _02896_
+ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__o21bai_1
XFILLER_195_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__03039_ _03039_ vssd1 vssd1 vccd1 vccd1 clknet_0__03039_ sky130_fd_sc_hd__clkbuf_16
XFILLER_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20291__306 clknet_1_1__leaf__03311_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__inv_2
X_21401_ net322 _01170_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1063 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21332_ net253 _01101_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_159_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21263_ clknet_leaf_88_i_clk _01032_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21194_ clknet_leaf_92_i_clk _00963_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_132_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ rbzero.tex_g0\[25\] rbzero.tex_g0\[24\] _03740_ vssd1 vssd1 vccd1 vccd1 _03744_
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ rbzero.tex_g0\[61\] rbzero.tex_g0\[60\] _04262_ vssd1 vssd1 vccd1 vccd1 _04558_
+ sky130_fd_sc_hd__mux2_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20978_ clknet_leaf_11_i_clk _00747_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10731_ _03707_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__clkbuf_1
XFILLER_198_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13450_ _06173_ _06186_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__xor2_1
X_10662_ _03671_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_201_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12401_ net34 _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__and2_1
XFILLER_22_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13381_ _06114_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__xnor2_2
X_10593_ _03634_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_166_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15120_ _07776_ _07777_ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__or2_1
X_12332_ net29 vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__inv_2
XFILLER_166_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15051_ _07713_ _07699_ _07698_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12263_ net21 vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__inv_2
XFILLER_126_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14002_ _06615_ _06738_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__or2_1
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ rbzero.wall_tracer.state\[8\] vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__inv_2
X_12194_ net18 net19 vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__nor2_1
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput62 net62 vssd1 vssd1 vccd1 vccd1 o_rgb[15] sky130_fd_sc_hd__buf_2
X_18810_ _02491_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__clkbuf_1
X_11145_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__inv_2
X_19790_ rbzero.pov.spi_buffer\[68\] rbzero.pov.spi_buffer\[69\] _03114_ vssd1 vssd1
+ vccd1 vccd1 _03124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18741_ _02428_ _02429_ _02430_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03290_ clknet_0__03290_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03290_
+ sky130_fd_sc_hd__clkbuf_16
X_11076_ _03888_ vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__clkbuf_1
X_15953_ _08590_ _08597_ vssd1 vssd1 vccd1 vccd1 _08598_ sky130_fd_sc_hd__xor2_1
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14904_ rbzero.wall_tracer.visualWallDist\[-6\] _07595_ vssd1 vssd1 vccd1 vccd1 _07611_
+ sky130_fd_sc_hd__or2_1
X_18672_ _08047_ _09565_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__nor2_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _08517_ _08525_ vssd1 vssd1 vccd1 vccd1 _08529_ sky130_fd_sc_hd__nor2_1
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ _10053_ _10056_ _10054_ vssd1 vssd1 vccd1 vccd1 _10188_ sky130_fd_sc_hd__a21boi_1
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ _07468_ _07557_ _07558_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__or3b_1
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ _10118_ _10114_ vssd1 vssd1 vccd1 vccd1 _10120_ sky130_fd_sc_hd__or2b_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14766_ _07473_ _07499_ _05814_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__a21oi_1
X_11978_ _04254_ _04748_ _04752_ _04371_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__a211o_1
XFILLER_189_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16505_ _09125_ _09148_ vssd1 vssd1 vccd1 vccd1 _09149_ sky130_fd_sc_hd__xnor2_2
XFILLER_189_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13717_ _06440_ _06452_ _06453_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10929_ _03811_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__clkbuf_1
X_17485_ _09958_ _09970_ vssd1 vssd1 vccd1 vccd1 _10051_ sky130_fd_sc_hd__nand2_1
X_14697_ _07394_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__nand2_1
XFILLER_147_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19224_ _02761_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16436_ _05397_ _05503_ _07971_ vssd1 vssd1 vccd1 vccd1 _09081_ sky130_fd_sc_hd__mux2_1
X_13648_ _06339_ _06383_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ rbzero.spi_registers.new_other\[10\] _02712_ vssd1 vssd1 vccd1 vccd1 _02718_
+ sky130_fd_sc_hd__or2_1
X_16367_ _07941_ _08097_ vssd1 vssd1 vccd1 vccd1 _09012_ sky130_fd_sc_hd__or2_1
X_13579_ _06309_ _06315_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__nand2_1
XFILLER_118_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_i_clk clknet_opt_12_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_173_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18106_ _01705_ _01714_ _01712_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a21o_1
XFILLER_145_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15318_ _07903_ rbzero.wall_tracer.stepDistY\[-6\] _05195_ vssd1 vssd1 vccd1 vccd1
+ _07963_ sky130_fd_sc_hd__a21o_1
X_19086_ _02675_ vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__clkbuf_1
X_16298_ _08811_ _08942_ vssd1 vssd1 vccd1 vccd1 _08943_ sky130_fd_sc_hd__xnor2_2
XFILLER_172_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18037_ _08242_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__buf_2
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15249_ _07894_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__buf_4
XFILLER_67_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_68_i_clk clknet_opt_11_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_i_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20134__165 clknet_1_0__leaf__03295_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__inv_2
XFILLER_114_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19988_ rbzero.pov.ready_buffer\[14\] _03252_ _03253_ rbzero.debug_overlay.vplaneX\[-6\]
+ _03254_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__o221a_1
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18939_ rbzero.pov.spi_buffer\[3\] rbzero.pov.ready_buffer\[3\] _02595_ vssd1 vssd1
+ vccd1 vccd1 _02599_ sky130_fd_sc_hd__mux2_1
XFILLER_140_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20901_ clknet_leaf_84_i_clk _00670_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.ready_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20832_ clknet_leaf_53_i_clk _00601_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistY\[-12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20763_ clknet_leaf_45_i_clk _00532_ vssd1 vssd1 vccd1 vccd1 rbzero.row_render.size\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20694_ clknet_leaf_58_i_clk _00478_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.stepDistX\[-1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21315_ net236 _01084_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21246_ clknet_leaf_79_i_clk _01015_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.facingY\[-9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_104_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21177_ clknet_leaf_5_i_clk _00946_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12950_ _05685_ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__xnor2_4
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11901_ _04675_ _04676_ _04139_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__mux2_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12881_ _05561_ _05461_ _05616_ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o22a_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _04306_ _04604_ _04608_ _04371_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a211o_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _05793_ _07356_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__and2_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14551_ _07080_ _07082_ _07084_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__o21a_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ rbzero.tex_g0\[17\] rbzero.tex_g0\[16\] _04129_ vssd1 vssd1 vccd1 vccd1 _04541_
+ sky130_fd_sc_hd__mux2_1
XFILLER_199_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _03698_ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__clkbuf_1
X_13502_ _06015_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__clkbuf_4
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14482_ _07164_ _07167_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__nand2_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ rbzero.wall_tracer.trackDistX\[-8\] _09844_ _05414_ vssd1 vssd1 vccd1 vccd1
+ _09845_ sky130_fd_sc_hd__mux2_1
XFILLER_186_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11694_ _04471_ _04463_ _04459_ rbzero.debug_overlay.vplaneY\[0\] _04472_ vssd1 vssd1
+ vccd1 vccd1 _04473_ sky130_fd_sc_hd__a221o_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_201_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16221_ _08860_ _08864_ vssd1 vssd1 vccd1 vccd1 _08866_ sky130_fd_sc_hd__nand2_1
X_13433_ _06168_ _06169_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__or2_1
X_10645_ _03662_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_195_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16152_ _08780_ _08781_ _08792_ _08794_ _08796_ vssd1 vssd1 vccd1 vccd1 _08797_ sky130_fd_sc_hd__a32oi_2
X_13364_ _05946_ _05961_ _06007_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__or3_1
X_10576_ rbzero.tex_r0\[3\] rbzero.tex_r0\[2\] _03624_ vssd1 vssd1 vccd1 vccd1 _03626_
+ sky130_fd_sc_hd__mux2_1
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12315_ net26 vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__clkbuf_4
X_15103_ _07758_ _07759_ _07760_ _07757_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__a22o_1
XFILLER_6_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16083_ _07958_ _08572_ vssd1 vssd1 vccd1 vccd1 _08728_ sky130_fd_sc_hd__or2_1
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13295_ _05978_ _06031_ _05962_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__o21bai_1
XFILLER_142_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15034_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__and2_1
X_19911_ rbzero.debug_overlay.playerY\[-3\] _03198_ _03211_ _03209_ vssd1 vssd1 vccd1
+ vccd1 _00995_ sky130_fd_sc_hd__o211a_1
X_12246_ _04977_ _05014_ _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__o21ai_1
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19842_ _07949_ _03143_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__nand2_1
X_12177_ _04908_ _04943_ _04947_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__a21oi_1
XFILLER_123_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ rbzero.wall_tracer.visualWallDist\[4\] rbzero.wall_tracer.visualWallDist\[3\]
+ rbzero.wall_tracer.visualWallDist\[2\] rbzero.wall_tracer.visualWallDist\[1\] vssd1
+ vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__or4_1
XFILLER_111_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19773_ _03115_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__clkbuf_1
X_16985_ _09620_ _09623_ vssd1 vssd1 vccd1 vccd1 _09625_ sky130_fd_sc_hd__or2_1
XFILLER_7_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18724_ _02407_ _02408_ _02409_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__o21bai_1
X_15936_ _08569_ _08577_ vssd1 vssd1 vccd1 vccd1 _08581_ sky130_fd_sc_hd__or2_1
XFILLER_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11059_ _03879_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18655_ _02139_ _02248_ _02140_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__o21a_1
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ _08460_ _08461_ vssd1 vssd1 vccd1 vccd1 _08512_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17606_ _05203_ _10171_ vssd1 vssd1 vccd1 vccd1 _10172_ sky130_fd_sc_hd__or2_1
XFILLER_36_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14818_ _05188_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__buf_4
X_18586_ _02269_ _02270_ _02281_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__and3_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_920 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15798_ _08259_ _08238_ vssd1 vssd1 vccd1 vccd1 _08443_ sky130_fd_sc_hd__nor2_1
XFILLER_205_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17537_ _10101_ _10102_ vssd1 vssd1 vccd1 vccd1 _10103_ sky130_fd_sc_hd__xor2_2
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14749_ _07468_ _07483_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__or2_1
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17468_ _05532_ _10033_ _10034_ _09817_ vssd1 vssd1 vccd1 vccd1 _10035_ sky130_fd_sc_hd__o31a_1
XFILLER_177_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19207_ rbzero.spi_registers.got_new_floor _02707_ vssd1 vssd1 vccd1 vccd1 _02751_
+ sky130_fd_sc_hd__nand2_2
XFILLER_73_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16419_ _09061_ _09062_ _09063_ vssd1 vssd1 vccd1 vccd1 _09064_ sky130_fd_sc_hd__and3_1
X_17399_ _08178_ _09103_ vssd1 vssd1 vccd1 vccd1 _09966_ sky130_fd_sc_hd__or2_1
XFILLER_164_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19138_ gpout0.vpos\[3\] _02704_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__and2_1
XFILLER_164_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19069_ rbzero.pov.spi_buffer\[65\] rbzero.pov.ready_buffer\[65\] _02660_ vssd1 vssd1
+ vccd1 vccd1 _02667_ sky130_fd_sc_hd__mux2_1
XFILLER_106_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_195_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21100_ net190 _00869_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b0\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21031_ clknet_leaf_11_i_clk _00800_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_vshift\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_102_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19586__42 clknet_1_1__leaf__03039_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__inv_2
XFILLER_43_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20815_ clknet_leaf_55_i_clk _00584_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.trackDistX\[-5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20746_ clknet_leaf_42_i_clk _00515_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.texu\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20677_ clknet_leaf_48_i_clk _00461_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.visualWallDist\[6\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__03293_ clknet_0__03293_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03293_
+ sky130_fd_sc_hd__clkbuf_16
X_10430_ rbzero.tex_r1\[5\] rbzero.tex_r1\[6\] _03538_ vssd1 vssd1 vccd1 vccd1 _03547_
+ sky130_fd_sc_hd__mux2_1
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10361_ rbzero.tex_r1\[38\] rbzero.tex_r1\[39\] _03505_ vssd1 vssd1 vccd1 vccd1 _03511_
+ sky130_fd_sc_hd__mux2_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12100_ gpout0.hpos\[3\] _04855_ _04857_ _04163_ vssd1 vssd1 vccd1 vccd1 _04872_
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ _05634_ _05775_ _05788_ _05789_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__or4_1
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12031_ rbzero.color_sky\[5\] rbzero.color_floor\[5\] _04144_ vssd1 vssd1 vccd1 vccd1
+ _04806_ sky130_fd_sc_hd__mux2_2
X_21229_ clknet_leaf_17_i_clk _00998_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.playerY\[0\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_104_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16770_ _09114_ _08178_ vssd1 vssd1 vccd1 vccd1 _09412_ sky130_fd_sc_hd__or2_1
XFILLER_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13982_ _06710_ _06713_ _06718_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__a21o_1
XFILLER_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20306__319 clknet_1_1__leaf__03313_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__inv_2
X_15721_ _08358_ _08365_ vssd1 vssd1 vccd1 vccd1 _08366_ sky130_fd_sc_hd__xnor2_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _05650_ _05669_ _05654_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__o21bai_1
XFILLER_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _02116_ _02117_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__or2_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15652_ _08281_ _08296_ vssd1 vssd1 vccd1 vccd1 _08297_ sky130_fd_sc_hd__xnor2_4
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _05577_ _05579_ _05582_ _05600_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__a211o_2
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _07206_ _07338_ _07339_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__o21ai_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _02068_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__xnor2_1
X_11815_ _04206_ _04592_ _04314_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a21o_1
XFILLER_15_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _08217_ _08225_ _08227_ vssd1 vssd1 vccd1 vccd1 _08228_ sky130_fd_sc_hd__o21a_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _05534_ _05536_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__nand2_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ rbzero.wall_tracer.trackDistX\[-2\] rbzero.wall_tracer.stepDistX\[-2\] vssd1
+ vssd1 vccd1 vccd1 _09891_ sky130_fd_sc_hd__and2_1
XFILLER_144_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14534_ _07268_ _07270_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__or2b_1
X_11746_ rbzero.tex_g0\[15\] _04135_ _04136_ _04126_ vssd1 vssd1 vccd1 vccd1 _04524_
+ sky130_fd_sc_hd__a31o_1
XFILLER_186_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17253_ _09829_ vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__clkbuf_1
X_11677_ rbzero.debug_overlay.vplaneX\[-6\] _04420_ _04447_ vssd1 vssd1 vccd1 vccd1
+ _04456_ sky130_fd_sc_hd__and3_1
X_14465_ _07147_ _07152_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__or2b_1
XFILLER_105_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16204_ _08778_ _08848_ vssd1 vssd1 vccd1 vccd1 _08849_ sky130_fd_sc_hd__xnor2_1
X_10628_ _03653_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__clkbuf_1
X_13416_ _05988_ _05980_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__nand2_4
XFILLER_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17184_ rbzero.traced_texa\[11\] _09770_ _09771_ rbzero.wall_tracer.visualWallDist\[11\]
+ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__a22o_1
X_14396_ _07129_ _07132_ _06239_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__a21oi_1
XFILLER_183_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16135_ _08743_ _08750_ vssd1 vssd1 vccd1 vccd1 _08780_ sky130_fd_sc_hd__nand2_1
X_13347_ _06059_ _06060_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__and2_1
X_10559_ rbzero.tex_r0\[11\] rbzero.tex_r0\[10\] _03613_ vssd1 vssd1 vccd1 vccd1 _03617_
+ sky130_fd_sc_hd__mux2_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13278_ _05750_ _05684_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__nor2_2
X_16066_ _08700_ _08709_ _08710_ vssd1 vssd1 vccd1 vccd1 _08711_ sky130_fd_sc_hd__a21o_1
XFILLER_115_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12229_ net44 _04963_ _04978_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__and3_1
X_15017_ _07680_ _07681_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__and2b_1
XFILLER_68_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19825_ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__buf_4
XFILLER_64_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19756_ _03106_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16968_ _09486_ _09495_ vssd1 vssd1 vccd1 vccd1 _09608_ sky130_fd_sc_hd__xnor2_1
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18707_ rbzero.wall_tracer.trackDistY\[-11\] rbzero.wall_tracer.stepDistY\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__or2_1
XFILLER_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15919_ _08492_ _08494_ vssd1 vssd1 vccd1 vccd1 _08564_ sky130_fd_sc_hd__nand2_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20246__266 clknet_1_1__leaf__03306_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__inv_2
X_19687_ _03047_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__clkbuf_4
XFILLER_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16899_ _08985_ _09420_ vssd1 vssd1 vccd1 vccd1 _09540_ sky130_fd_sc_hd__and2_1
X_18638_ _09141_ _08423_ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__nor2_1
XFILLER_37_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18569_ _02071_ _02172_ _02174_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a21bo_1
XFILLER_33_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20600_ gpout2.clk_div\[0\] net60 vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__nor2_1
XFILLER_21_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21580_ net501 _01349_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20531_ rbzero.texV\[7\] _03327_ _03332_ _03423_ vssd1 vssd1 vccd1 vccd1 _01403_
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20462_ _03362_ _03363_ _03364_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__o21ai_1
XFILLER_181_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_4_0_i_clk clknet_3_2_0_i_clk vssd1 vssd1 vccd1 vccd1 clknet_opt_4_0_i_clk
+ sky130_fd_sc_hd__clkbuf_16
X_20393_ clknet_1_0__leaf__04835_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__buf_1
XFILLER_145_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21014_ clknet_leaf_8_i_clk _00783_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.new_leak\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11600_ _04224_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__buf_4
XFILLER_54_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ _05322_ _05332_ _05320_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a21oi_1
XFILLER_168_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11531_ _04206_ _04270_ _04310_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nand3b_1
XFILLER_141_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20729_ clknet_leaf_84_i_clk _00498_ vssd1 vssd1 vccd1 vccd1 rbzero.wall_tracer.rayAddendX\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14250_ _06953_ _06959_ _06958_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__a21o_1
X_11462_ _04241_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__buf_4
XFILLER_104_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13201_ _05925_ _05927_ _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__a21bo_1
XFILLER_183_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10413_ _03482_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__clkbuf_4
X_14181_ _06704_ _06672_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__nor2_1
XFILLER_164_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11393_ gpout0.hpos\[7\] _04159_ _04171_ _04172_ vssd1 vssd1 vccd1 vccd1 _04173_
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13132_ _05820_ _05868_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__nand2_1
X_10344_ rbzero.tex_r1\[46\] rbzero.tex_r1\[47\] _03494_ vssd1 vssd1 vccd1 vccd1 _03502_
+ sky130_fd_sc_hd__mux2_1
XFILLER_164_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17940_ _01634_ _01641_ _01642_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__nand3_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__buf_4
XFILLER_151_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12014_ rbzero.tex_b1\[41\] rbzero.tex_b1\[40\] _04392_ vssd1 vssd1 vccd1 vccd1 _04789_
+ sky130_fd_sc_hd__mux2_1
X_17871_ _01496_ _01511_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__nor2_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16822_ _09335_ _09337_ _09334_ vssd1 vssd1 vccd1 vccd1 _09464_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19541_ _02906_ _03014_ _03015_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__mux2_1
X_16753_ _08383_ _08570_ vssd1 vssd1 vccd1 vccd1 _09395_ sky130_fd_sc_hd__nor2_1
XFILLER_115_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13965_ _06700_ _06701_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__nand2_1
XFILLER_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_207_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15704_ _08337_ _08347_ _08348_ vssd1 vssd1 vccd1 vccd1 _08349_ sky130_fd_sc_hd__a21o_1
XFILLER_19_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__03041_ clknet_0__03041_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03041_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19472_ _02950_ _02951_ _02952_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__nand3_1
X_12916_ rbzero.wall_tracer.visualWallDist\[7\] _05571_ _05572_ vssd1 vssd1 vccd1
+ vccd1 _05653_ sky130_fd_sc_hd__a21o_1
X_16684_ _09324_ _09326_ vssd1 vssd1 vccd1 vccd1 _09327_ sky130_fd_sc_hd__xor2_1
X_13896_ _06620_ _06631_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__nand2_1
XFILLER_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18423_ _02120_ _02121_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__nand2_1
XFILLER_206_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15635_ _08262_ _08278_ _08279_ vssd1 vssd1 vccd1 vccd1 _08280_ sky130_fd_sc_hd__a21oi_2
XFILLER_34_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12847_ _05475_ _05583_ _05561_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__mux2_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18354_ _02044_ _02052_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__xor2_1
XFILLER_199_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ _07894_ _05454_ vssd1 vssd1 vccd1 vccd1 _08211_ sky130_fd_sc_hd__nand2_1
XFILLER_187_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ rbzero.debug_overlay.playerX\[4\] _05522_ _05394_ vssd1 vssd1 vccd1 vccd1
+ _05523_ sky130_fd_sc_hd__mux2_1
XFILLER_203_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19580__37 clknet_1_0__leaf__03038_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__inv_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _09874_ _09875_ vssd1 vssd1 vccd1 vccd1 _09876_ sky130_fd_sc_hd__xnor2_1
X_14517_ _07060_ _06843_ _07066_ _07253_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__a31o_1
XFILLER_202_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18285_ _01860_ _01620_ _01984_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__or3_1
XFILLER_148_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11729_ rbzero.debug_overlay.playerY\[-6\] _04475_ _04498_ _04507_ vssd1 vssd1 vccd1
+ vccd1 _04508_ sky130_fd_sc_hd__a211o_1
XFILLER_187_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15497_ _08113_ _08139_ _08140_ _08141_ vssd1 vssd1 vccd1 vccd1 _08142_ sky130_fd_sc_hd__o22a_1
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17236_ rbzero.wall_tracer.trackDistX\[-11\] rbzero.wall_tracer.stepDistX\[-11\]
+ vssd1 vssd1 vccd1 vccd1 _09814_ sky130_fd_sc_hd__nand2_1
XFILLER_31_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14448_ _07112_ _07113_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__and2_1
XFILLER_174_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17167_ rbzero.traced_texa\[-3\] _09768_ _09767_ rbzero.wall_tracer.visualWallDist\[-3\]
+ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__a22o_1
XFILLER_122_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14379_ _06698_ _07072_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__nor2_1
XFILLER_116_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16118_ _08737_ _08761_ _08762_ vssd1 vssd1 vccd1 vccd1 _08763_ sky130_fd_sc_hd__a21oi_2
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17098_ _09594_ _09596_ _09592_ vssd1 vssd1 vccd1 vccd1 _09738_ sky130_fd_sc_hd__a21oi_2
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16049_ _08682_ _08689_ _08691_ vssd1 vssd1 vccd1 vccd1 _08694_ sky130_fd_sc_hd__and3_1
XFILLER_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19808_ net52 rbzero.pov.sclk_buffer\[0\] _02695_ vssd1 vssd1 vccd1 vccd1 _03133_
+ sky130_fd_sc_hd__mux2_1
XFILLER_97_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__03308_ clknet_0__03308_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__03308_
+ sky130_fd_sc_hd__clkbuf_16
X_19739_ _03097_ vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_53_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21632_ clknet_leaf_30_i_clk _01401_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_178_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21563_ net484 _01332_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r1\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20514_ _03406_ _03409_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__xnor2_1
X_21494_ net415 _01263_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20445_ rbzero.traced_texa\[-6\] rbzero.texV\[-6\] vssd1 vssd1 vccd1 vccd1 _03351_
+ sky130_fd_sc_hd__nor2_1
XFILLER_147_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20229__250 clknet_1_1__leaf__03305_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__inv_2
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13750_ _06468_ _06482_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__xor2_1
XFILLER_84_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10962_ rbzero.tex_b1\[11\] rbzero.tex_b1\[12\] _03828_ vssd1 vssd1 vccd1 vccd1 _03829_
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ rbzero.debug_overlay.facingX\[10\] _05448_ vssd1 vssd1 vccd1 vccd1 _05449_
+ sky130_fd_sc_hd__nand2_1
XFILLER_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13681_ _06394_ _06416_ _06417_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__o21a_1
X_10893_ _03792_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_203_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15420_ rbzero.debug_overlay.playerX\[-3\] _07946_ vssd1 vssd1 vccd1 vccd1 _08065_
+ sky130_fd_sc_hd__nand2_1
X_12632_ _05383_ _05384_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__xnor2_1
XFILLER_58_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_203_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15351_ _07995_ vssd1 vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12563_ _05315_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__or2_1
XFILLER_129_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11514_ _04292_ _04293_ _04266_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__mux2_1
XFILLER_157_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14302_ _07036_ _07037_ _06882_ _07034_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__a211o_1
X_18070_ _01632_ _01651_ _01650_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__a21o_1
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15282_ _07541_ _07926_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1 _07927_
+ sky130_fd_sc_hd__mux2_1
X_12494_ rbzero.wall_tracer.trackDistY\[-6\] _05237_ rbzero.wall_tracer.trackDistY\[-7\]
+ _05238_ _05248_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a221o_1
XFILLER_102_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17021_ _07976_ vssd1 vssd1 vccd1 vccd1 _09661_ sky130_fd_sc_hd__clkbuf_4
X_11445_ _04224_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__buf_4
X_14233_ _06944_ _06969_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__nand2_1
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14164_ _06892_ _06899_ _06900_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__a21oi_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11376_ rbzero.row_render.size\[8\] rbzero.row_render.size\[7\] rbzero.row_render.size\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__nand3_1
XFILLER_98_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10327_ rbzero.tex_r1\[54\] rbzero.tex_r1\[55\] _03483_ vssd1 vssd1 vccd1 vccd1 _03493_
+ sky130_fd_sc_hd__mux2_1
X_13115_ _05847_ _05848_ _05851_ _05700_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__a211o_2
XFILLER_180_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14095_ _06826_ _06831_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__xor2_1
X_18972_ _02594_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__clkbuf_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17923_ _01624_ _01625_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__xnor2_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _05711_ _05712_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__xnor2_2
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17854_ _01556_ _01557_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__xnor2_1
XFILLER_26_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16805_ _09445_ _09446_ vssd1 vssd1 vccd1 vccd1 _09447_ sky130_fd_sc_hd__xor2_1
XFILLER_66_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17785_ _01487_ _01488_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__nor2_1
X_14997_ rbzero.wall_tracer.stepDistX\[5\] _07568_ _07660_ vssd1 vssd1 vccd1 vccd1
+ _07669_ sky130_fd_sc_hd__mux2_1
XFILLER_35_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19524_ rbzero.wall_tracer.rayAddendY\[8\] rbzero.wall_tracer.rayAddendY\[7\] _02906_
+ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__o21ai_1
X_16736_ _09362_ _09377_ vssd1 vssd1 vccd1 vccd1 _09378_ sky130_fd_sc_hd__xnor2_1
X_13948_ _06665_ _06670_ _06684_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__a21o_1
XFILLER_47_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19455_ _02923_ _02925_ _02935_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16667_ _09305_ _09306_ _09308_ vssd1 vssd1 vccd1 vccd1 _09310_ sky130_fd_sc_hd__a21o_1
X_13879_ _06273_ _06593_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__nand2_1
XFILLER_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18406_ _02102_ _02104_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__xor2_2
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15618_ rbzero.debug_overlay.playerX\[-9\] _08147_ _07979_ vssd1 vssd1 vccd1 vccd1
+ _08263_ sky130_fd_sc_hd__a21o_2
XFILLER_195_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19386_ rbzero.debug_overlay.vplaneY\[-5\] rbzero.debug_overlay.vplaneY\[-9\] vssd1
+ vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__or2_1
X_16598_ _09118_ _09123_ vssd1 vssd1 vccd1 vccd1 _09241_ sky130_fd_sc_hd__nand2_1
X_18337_ _01756_ _01970_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__nand2_1
XFILLER_175_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20358__367 clknet_1_1__leaf__03317_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__inv_2
X_15549_ _08008_ vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__buf_4
XFILLER_33_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18268_ _01879_ _01880_ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__a21bo_1
XFILLER_148_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17219_ _09779_ _09798_ _09799_ _09781_ rbzero.wall_tracer.mapX\[10\] vssd1 vssd1
+ vccd1 vccd1 _00575_ sky130_fd_sc_hd__a32o_1
XFILLER_162_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18199_ _01897_ _01899_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__xnor2_1
XFILLER_190_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_196_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20161_ clknet_1_1__leaf__03298_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__buf_1
XFILLER_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20387__13 clknet_1_1__leaf__03320_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__inv_2
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994_ clknet_leaf_13_i_clk _00763_ vssd1 vssd1 vccd1 vccd1 rbzero.spi_registers.vshift\[5\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_198_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21615_ clknet_leaf_27_i_clk _01384_ vssd1 vssd1 vccd1 vccd1 rbzero.texV\[-12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21546_ net467 _01315_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_194_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21477_ net398 _01246_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g1\[56\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11230_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__buf_6
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20428_ rbzero.texV\[-10\] _03175_ _03332_ _03337_ vssd1 vssd1 vccd1 vccd1 _01386_
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__03044_ clknet_0__03044_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__03044_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_136_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11161_ rbzero.wall_tracer.mapY\[9\] rbzero.wall_tracer.mapY\[8\] rbzero.wall_tracer.mapY\[11\]
+ rbzero.wall_tracer.mapY\[10\] vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__or4_1
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11092_ _03896_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_1_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14920_ rbzero.wall_tracer.visualWallDist\[-2\] _07618_ vssd1 vssd1 vccd1 vccd1 _07623_
+ sky130_fd_sc_hd__or2_1
XFILLER_49_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14851_ _05742_ _07383_ _07390_ _05736_ _05737_ vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__a2111oi_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13802_ _06406_ _06531_ _06530_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__nand3b_1
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ _10133_ _10135_ vssd1 vssd1 vccd1 vccd1 _10136_ sky130_fd_sc_hd__and2_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14782_ rbzero.wall_tracer.stepDistY\[-8\] _00004_ vssd1 vssd1 vccd1 vccd1 _07515_
+ sky130_fd_sc_hd__nor2_1
X_11994_ _04766_ _04767_ _04768_ _04225_ _04229_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__o221a_1
XFILLER_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16521_ _09164_ vssd1 vssd1 vccd1 vccd1 _09165_ sky130_fd_sc_hd__clkbuf_4
X_13733_ _06057_ _06031_ _05945_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__o21ai_1
XFILLER_182_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10945_ rbzero.tex_b1\[19\] rbzero.tex_b1\[20\] _03817_ vssd1 vssd1 vccd1 vccd1 _03820_
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19240_ _02771_ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__clkbuf_1
X_16452_ _08821_ vssd1 vssd1 vccd1 vccd1 _09096_ sky130_fd_sc_hd__clkbuf_4
XFILLER_32_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13664_ _05990_ _06009_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__or2_1
XFILLER_182_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10876_ _03783_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15403_ _07486_ _07455_ _07483_ rbzero.wall_tracer.state\[3\] vssd1 vssd1 vccd1 vccd1
+ _08048_ sky130_fd_sc_hd__a211oi_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _05367_ _05368_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__nand2_1
X_19171_ _02727_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__buf_4
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16383_ _08147_ _09027_ vssd1 vssd1 vccd1 vccd1 _09028_ sky130_fd_sc_hd__or2_2
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _06148_ _06147_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__xnor2_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18122_ _01462_ _09526_ _09621_ rbzero.wall_tracer.visualWallDist\[10\] vssd1 vssd1
+ vccd1 vccd1 _01823_ sky130_fd_sc_hd__and4bb_1
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15334_ rbzero.debug_overlay.playerY\[-9\] _04013_ _05196_ _07978_ vssd1 vssd1 vccd1
+ vccd1 _07979_ sky130_fd_sc_hd__o211a_1
X_12546_ _05296_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__and2_1
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18053_ _01636_ _01639_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__nand2_1
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15265_ _07904_ _07909_ vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__nand2_1
X_12477_ _05216_ _05229_ _05231_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__o21a_1
XFILLER_138_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17004_ _09642_ _09643_ vssd1 vssd1 vccd1 vccd1 _09644_ sky130_fd_sc_hd__and2b_1
XANTENNA_4 _05533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _06951_ _06952_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__nor2_1
XFILLER_32_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11428_ _04141_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__buf_6
X_15196_ _07847_ _07848_ _07833_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__o21bai_1
XFILLER_99_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14147_ _06856_ _06879_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__xnor2_1
XFILLER_98_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11359_ _04138_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__buf_6
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14078_ _06813_ _06800_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__or2b_1
X_18955_ _02607_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17906_ _01573_ _01608_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__nand2_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13029_ _05765_ _05576_ _05657_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__o21ba_1
X_18886_ _02556_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17837_ _10233_ _10280_ _01540_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__a21boi_1
XFILLER_67_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17768_ _10074_ _10217_ _10219_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__o21ai_1
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16719_ _09358_ _09360_ vssd1 vssd1 vccd1 vccd1 _09361_ sky130_fd_sc_hd__xor2_1
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19507_ _02984_ _02985_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__nand2_1
XFILLER_81_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17699_ _10257_ _10263_ vssd1 vssd1 vccd1 vccd1 _10264_ sky130_fd_sc_hd__xor2_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19438_ rbzero.wall_tracer.rayAddendY\[2\] rbzero.wall_tracer.rayAddendY\[1\] rbzero.debug_overlay.vplaneY\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__o21ai_1
XFILLER_90_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__03038_ _03038_ vssd1 vssd1 vccd1 vccd1 clknet_0__03038_ sky130_fd_sc_hd__clkbuf_16
X_19369_ _07676_ _02849_ _02850_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a31o_1
XFILLER_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21400_ net321 _01169_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_g0\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21331_ net252 _01100_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_b1\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_190_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_194_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21262_ clknet_leaf_96_i_clk _01031_ vssd1 vssd1 vccd1 vccd1 rbzero.debug_overlay.vplaneX\[-4\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_163_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21193_ clknet_leaf_78_i_clk _00962_ vssd1 vssd1 vccd1 vccd1 rbzero.pov.spi_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20111__144 clknet_1_0__leaf__03293_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__inv_2
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ clknet_leaf_10_i_clk _00746_ vssd1 vssd1 vccd1 vccd1 rbzero.color_sky\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10730_ rbzero.tex_g0\[58\] rbzero.tex_g0\[57\] _03706_ vssd1 vssd1 vccd1 vccd1 _03707_
+ sky130_fd_sc_hd__mux2_1
XFILLER_207_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10661_ rbzero.tex_g1\[26\] rbzero.tex_g1\[27\] _03669_ vssd1 vssd1 vccd1 vccd1 _03671_
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12400_ _04154_ _03477_ _05143_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__mux2_1
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13380_ _06115_ _05923_ _06116_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__and3_1
X_10592_ rbzero.tex_g1\[58\] rbzero.tex_g1\[59\] _03549_ vssd1 vssd1 vccd1 vccd1 _03634_
+ sky130_fd_sc_hd__mux2_1
XFILLER_103_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ _05082_ _05087_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__nand2_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21529_ net450 _01298_ vssd1 vssd1 vccd1 vccd1 rbzero.tex_r0\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12262_ net23 _05023_ _05026_ _05030_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__o211a_1
XFILLER_5_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15050_ rbzero.debug_overlay.vplaneX\[-4\] rbzero.wall_tracer.rayAddendX\[-4\] vssd1
+ vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__or2_1
XFILLER_182_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14001_ _06614_ _06598_ _06599_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__and3_1
X_11213_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__clkbuf_4
X_12193_ net17 net16 vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__nor2_1
XFILLER_134_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11144_ rbzero.map_rom.b6 vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__clkbuf_4
Xoutput63 net63 vssd1 vssd1 vccd1 vccd1 o_rgb[22] sky130_fd_sc_hd__buf_2
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18740_ _02421_ _02423_ _02422_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__o21bai_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11075_ rbzero.tex_b0\[22\] rbzero.tex_b0\[21\] _03887_ vssd1 vssd1 vccd1 vccd1 _03888_
+ sky130_fd_sc_hd__mux2_1
X_15952_ _08593_ _08595_ _08596_ vssd1 vssd1 vccd1 vccd1 _08597_ sky130_fd_sc_hd__o21a_1
XFILLER_23_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14903_ rbzero.wall_tracer.trackDistY\[-6\] rbzero.wall_tracer.trackDistX\[-6\] _07592_
+ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__mux2_1
X_20086__121 clknet_1_1__leaf__03291_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__inv_2
X_18671_ _02144_ _02366_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__xnor2_1
XFILLER_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _08527_ _08474_ vssd1 vssd1 vccd1 vccd1 _08528_ sky130_fd_sc_hd__xnor2_2
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17622_ _10087_ _10050_ vssd1 vssd1 vccd1 vccd1 _10187_ sky130_fd_sc_hd__or2b_1
XFILLER_64_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14834_ _05834_ _05800_ _07520_ vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__or3_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17553_ _10114_ _10118_ vssd1 vssd1 vccd1 vccd1 _10119_ sky130_fd_sc_hd__and2b_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _07497_ _07498_ _05952_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__mux2_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11977_ _04225_ _04749_ _04750_ _04751_ _04208_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__o221a_1
XFILLER_189_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16504_ _09145_ _09147_ vssd1 vssd1 vccd1 vccd1 _09148_ sky130_fd_sc_hd__xor2_2
XFILLER_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13716_ _06441_ _06451_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__and2_1
XFILLER_204_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17484_ _09938_ _09950_ _10049_ vssd1 vssd1 vccd1 vccd1 _10050_ sky130_fd_sc_hd__a21o_1
X_10928_ rbzero.tex_b1\[27\] rbzero.tex_b1\[28\] _03806_ vssd1 vssd1 vccd1 vccd1 _03811_
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14696_ _07375_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__clkbuf_4
XFILLER_189_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19223_ rbzero.spi_registers.got_new_vshift _02708_ vssd1 vssd1 vccd1 vccd1 _02761_
+ sky130_fd_sc_hd__and2_1
XFILLER_149_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16435_ _09066_ _09079_ vssd1 vssd1 vccd1 vccd1 _09080_ sky130_fd_sc_hd__xor2_2
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13647_ _05824_ _05940_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__or2_1
XFILLER_32_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10859_ rbzero.tex_b1\[60\] rbzero.tex_b1\[61\] _03773_ vssd1 vssd1 vccd1 vccd1 _03775_
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19154_ rbzero.otherx\[3\] _02710_ _02717_ _02714_ vssd1 vssd1 vccd1 vccd1 _00732_
+ sky130_fd_sc_hd__o211a_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _08360_ _09009_ _09010_ vssd1 vssd1 vccd1 vccd1 _09011_ sky130_fd_sc_hd__a21o_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _06101_ _06310_ _06311_ _06314_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__o22a_1
XFILLER_185_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18105_ _01698_ _01732_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__nand2_1
XFILLER_9_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15317_ _07933_ _07530_ _07961_ vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__o21ai_4
XFILLER_172_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19085_ rbzero.pov.spi_buffer\[73\] rbzero.pov.ready_buffer\[73\] _02594_ vssd1 vssd1
+ vccd1 vccd1 _02675_ sky130_fd_sc_hd__mux2_1
X_12529_ _05283_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__clkbuf_4
X_16297_ _08764_ _08807_ _08941_ vssd1 vssd1 vccd1 vccd1 _08942_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18036_ _08242_ _01737_ _10238_ _09552_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__or4_1
XFILLER_145_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15248_ _07893_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__clkbuf_4
XFILLER_132_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15179_ _07820_ rbzero.debug_overlay.vplaneX\[-2\] vssd1 vssd1 vccd1 vccd1 _07833_
+ sky130_fd_sc_hd__nor2_1
XFILLER_158_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19987_ rbzero.pov.ready_buffer\[13\] _03252_ _03253_ rbzero.debug_overlay.vplaneX\[-7\]
+ _03254_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__o221a_1
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18938_ _02598_ vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__clkbuf_1
.ends


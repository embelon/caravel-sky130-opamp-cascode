VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_io_control
  CLASS BLOCK ;
  FOREIGN analog_io_control ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 240.000 ;
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 34.040 80.000 34.640 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 72.120 80.000 72.720 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 110.200 80.000 110.800 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 148.280 80.000 148.880 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 186.360 80.000 186.960 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 224.440 80.000 225.040 ;
    END
  END io_oeb[5]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 15.000 80.000 15.600 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 53.080 80.000 53.680 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 91.160 80.000 91.760 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 129.240 80.000 129.840 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 167.320 80.000 167.920 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 205.400 80.000 206.000 ;
    END
  END io_out[5]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 13.285 10.640 14.885 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 30.420 10.640 32.020 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.555 10.640 49.155 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.690 10.640 66.290 228.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.850 10.640 23.450 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.985 10.640 40.585 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.120 10.640 57.720 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.255 10.640 74.855 228.720 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 224.345 74.250 227.175 ;
        RECT 5.330 218.905 74.250 221.735 ;
        RECT 5.330 213.465 74.250 216.295 ;
        RECT 5.330 208.025 74.250 210.855 ;
        RECT 5.330 202.585 74.250 205.415 ;
        RECT 5.330 197.145 74.250 199.975 ;
        RECT 5.330 191.705 74.250 194.535 ;
        RECT 5.330 186.265 74.250 189.095 ;
        RECT 5.330 180.825 74.250 183.655 ;
        RECT 5.330 175.385 74.250 178.215 ;
        RECT 5.330 169.945 74.250 172.775 ;
        RECT 5.330 164.505 74.250 167.335 ;
        RECT 5.330 159.065 74.250 161.895 ;
        RECT 5.330 153.625 74.250 156.455 ;
        RECT 5.330 148.185 74.250 151.015 ;
        RECT 5.330 142.745 74.250 145.575 ;
        RECT 5.330 137.305 74.250 140.135 ;
        RECT 5.330 131.865 74.250 134.695 ;
        RECT 5.330 126.425 74.250 129.255 ;
        RECT 5.330 120.985 74.250 123.815 ;
        RECT 5.330 115.545 74.250 118.375 ;
        RECT 5.330 110.105 74.250 112.935 ;
        RECT 5.330 104.665 74.250 107.495 ;
        RECT 5.330 99.225 74.250 102.055 ;
        RECT 5.330 93.785 74.250 96.615 ;
        RECT 5.330 88.345 74.250 91.175 ;
        RECT 5.330 82.905 74.250 85.735 ;
        RECT 5.330 77.465 74.250 80.295 ;
        RECT 5.330 72.025 74.250 74.855 ;
        RECT 5.330 66.585 74.250 69.415 ;
        RECT 5.330 61.145 74.250 63.975 ;
        RECT 5.330 55.705 74.250 58.535 ;
        RECT 5.330 50.265 74.250 53.095 ;
        RECT 5.330 44.825 74.250 47.655 ;
        RECT 5.330 39.385 74.250 42.215 ;
        RECT 5.330 33.945 74.250 36.775 ;
        RECT 5.330 28.505 74.250 31.335 ;
        RECT 5.330 23.065 74.250 25.895 ;
        RECT 5.330 17.625 74.250 20.455 ;
        RECT 5.330 12.185 74.250 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 74.060 228.565 ;
      LAYER met1 ;
        RECT 5.520 10.640 74.855 228.720 ;
      LAYER met2 ;
        RECT 13.315 10.695 74.825 228.665 ;
      LAYER met3 ;
        RECT 13.295 225.440 76.000 228.645 ;
        RECT 13.295 224.040 75.600 225.440 ;
        RECT 13.295 206.400 76.000 224.040 ;
        RECT 13.295 205.000 75.600 206.400 ;
        RECT 13.295 187.360 76.000 205.000 ;
        RECT 13.295 185.960 75.600 187.360 ;
        RECT 13.295 168.320 76.000 185.960 ;
        RECT 13.295 166.920 75.600 168.320 ;
        RECT 13.295 149.280 76.000 166.920 ;
        RECT 13.295 147.880 75.600 149.280 ;
        RECT 13.295 130.240 76.000 147.880 ;
        RECT 13.295 128.840 75.600 130.240 ;
        RECT 13.295 111.200 76.000 128.840 ;
        RECT 13.295 109.800 75.600 111.200 ;
        RECT 13.295 92.160 76.000 109.800 ;
        RECT 13.295 90.760 75.600 92.160 ;
        RECT 13.295 73.120 76.000 90.760 ;
        RECT 13.295 71.720 75.600 73.120 ;
        RECT 13.295 54.080 76.000 71.720 ;
        RECT 13.295 52.680 75.600 54.080 ;
        RECT 13.295 35.040 76.000 52.680 ;
        RECT 13.295 33.640 75.600 35.040 ;
        RECT 13.295 16.000 76.000 33.640 ;
        RECT 13.295 14.600 75.600 16.000 ;
        RECT 13.295 10.715 76.000 14.600 ;
  END
END analog_io_control
END LIBRARY


// This is the unpowered netlist.
module top_ew_algofoogle (i_clk,
    i_debug_map_overlay,
    i_debug_trace_overlay,
    i_debug_vec_overlay,
    i_la_invalid,
    i_reg_csb,
    i_reg_mosi,
    i_reg_outs_enb,
    i_reg_sclk,
    i_reset_lock_a,
    i_reset_lock_b,
    i_spare_0,
    i_spare_1,
    i_vec_csb,
    i_vec_mosi,
    i_vec_sclk,
    o_hsync,
    o_reset,
    o_tex_csb,
    o_tex_oeb0,
    o_tex_out0,
    o_tex_sclk,
    o_vsync,
    i_gpout0_sel,
    i_gpout1_sel,
    i_gpout2_sel,
    i_gpout3_sel,
    i_gpout4_sel,
    i_gpout5_sel,
    i_mode,
    i_tex_in,
    o_gpout,
    o_rgb,
    ones,
    zeros);
 input i_clk;
 input i_debug_map_overlay;
 input i_debug_trace_overlay;
 input i_debug_vec_overlay;
 input i_la_invalid;
 input i_reg_csb;
 input i_reg_mosi;
 input i_reg_outs_enb;
 input i_reg_sclk;
 input i_reset_lock_a;
 input i_reset_lock_b;
 input i_spare_0;
 input i_spare_1;
 input i_vec_csb;
 input i_vec_mosi;
 input i_vec_sclk;
 output o_hsync;
 output o_reset;
 output o_tex_csb;
 output o_tex_oeb0;
 output o_tex_out0;
 output o_tex_sclk;
 output o_vsync;
 input [5:0] i_gpout0_sel;
 input [5:0] i_gpout1_sel;
 input [5:0] i_gpout2_sel;
 input [5:0] i_gpout3_sel;
 input [5:0] i_gpout4_sel;
 input [5:0] i_gpout5_sel;
 input [2:0] i_mode;
 input [3:0] i_tex_in;
 output [5:0] o_gpout;
 output [23:0] o_rgb;
 output [15:0] ones;
 output [15:0] zeros;

 wire _00000_;
 wire _00001_;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire clknet_leaf_0_i_clk;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire \gpout0.clk_div[0] ;
 wire \gpout0.clk_div[1] ;
 wire \gpout0.hpos[0] ;
 wire \gpout0.hpos[1] ;
 wire \gpout0.hpos[2] ;
 wire \gpout0.hpos[3] ;
 wire \gpout0.hpos[4] ;
 wire \gpout0.hpos[5] ;
 wire \gpout0.hpos[6] ;
 wire \gpout0.hpos[7] ;
 wire \gpout0.hpos[8] ;
 wire \gpout0.hpos[9] ;
 wire \gpout0.vpos[0] ;
 wire \gpout0.vpos[1] ;
 wire \gpout0.vpos[2] ;
 wire \gpout0.vpos[3] ;
 wire \gpout0.vpos[4] ;
 wire \gpout0.vpos[5] ;
 wire \gpout0.vpos[6] ;
 wire \gpout0.vpos[7] ;
 wire \gpout0.vpos[8] ;
 wire \gpout0.vpos[9] ;
 wire \gpout1.clk_div[0] ;
 wire \gpout1.clk_div[1] ;
 wire \gpout2.clk_div[0] ;
 wire \gpout2.clk_div[1] ;
 wire \gpout3.clk_div[0] ;
 wire \gpout3.clk_div[1] ;
 wire \gpout4.clk_div[0] ;
 wire \gpout4.clk_div[1] ;
 wire \gpout5.clk_div[0] ;
 wire \gpout5.clk_div[1] ;
 wire net76;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net77;
 wire net92;
 wire net93;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net110;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire \rbzero.color_floor[0] ;
 wire \rbzero.color_floor[1] ;
 wire \rbzero.color_floor[2] ;
 wire \rbzero.color_floor[3] ;
 wire \rbzero.color_floor[4] ;
 wire \rbzero.color_floor[5] ;
 wire \rbzero.color_sky[0] ;
 wire \rbzero.color_sky[1] ;
 wire \rbzero.color_sky[2] ;
 wire \rbzero.color_sky[3] ;
 wire \rbzero.color_sky[4] ;
 wire \rbzero.color_sky[5] ;
 wire \rbzero.debug_overlay.facingX[-1] ;
 wire \rbzero.debug_overlay.facingX[-2] ;
 wire \rbzero.debug_overlay.facingX[-3] ;
 wire \rbzero.debug_overlay.facingX[-4] ;
 wire \rbzero.debug_overlay.facingX[-5] ;
 wire \rbzero.debug_overlay.facingX[-6] ;
 wire \rbzero.debug_overlay.facingX[-7] ;
 wire \rbzero.debug_overlay.facingX[-8] ;
 wire \rbzero.debug_overlay.facingX[-9] ;
 wire \rbzero.debug_overlay.facingX[0] ;
 wire \rbzero.debug_overlay.facingX[10] ;
 wire \rbzero.debug_overlay.facingY[-1] ;
 wire \rbzero.debug_overlay.facingY[-2] ;
 wire \rbzero.debug_overlay.facingY[-3] ;
 wire \rbzero.debug_overlay.facingY[-4] ;
 wire \rbzero.debug_overlay.facingY[-5] ;
 wire \rbzero.debug_overlay.facingY[-6] ;
 wire \rbzero.debug_overlay.facingY[-7] ;
 wire \rbzero.debug_overlay.facingY[-8] ;
 wire \rbzero.debug_overlay.facingY[-9] ;
 wire \rbzero.debug_overlay.facingY[0] ;
 wire \rbzero.debug_overlay.facingY[10] ;
 wire \rbzero.debug_overlay.playerX[-1] ;
 wire \rbzero.debug_overlay.playerX[-2] ;
 wire \rbzero.debug_overlay.playerX[-3] ;
 wire \rbzero.debug_overlay.playerX[-4] ;
 wire \rbzero.debug_overlay.playerX[-5] ;
 wire \rbzero.debug_overlay.playerX[-6] ;
 wire \rbzero.debug_overlay.playerX[-7] ;
 wire \rbzero.debug_overlay.playerX[-8] ;
 wire \rbzero.debug_overlay.playerX[-9] ;
 wire \rbzero.debug_overlay.playerX[0] ;
 wire \rbzero.debug_overlay.playerX[1] ;
 wire \rbzero.debug_overlay.playerX[2] ;
 wire \rbzero.debug_overlay.playerX[3] ;
 wire \rbzero.debug_overlay.playerX[4] ;
 wire \rbzero.debug_overlay.playerX[5] ;
 wire \rbzero.debug_overlay.playerY[-1] ;
 wire \rbzero.debug_overlay.playerY[-2] ;
 wire \rbzero.debug_overlay.playerY[-3] ;
 wire \rbzero.debug_overlay.playerY[-4] ;
 wire \rbzero.debug_overlay.playerY[-5] ;
 wire \rbzero.debug_overlay.playerY[-6] ;
 wire \rbzero.debug_overlay.playerY[-7] ;
 wire \rbzero.debug_overlay.playerY[-8] ;
 wire \rbzero.debug_overlay.playerY[-9] ;
 wire \rbzero.debug_overlay.playerY[0] ;
 wire \rbzero.debug_overlay.playerY[1] ;
 wire \rbzero.debug_overlay.playerY[2] ;
 wire \rbzero.debug_overlay.playerY[3] ;
 wire \rbzero.debug_overlay.playerY[4] ;
 wire \rbzero.debug_overlay.playerY[5] ;
 wire \rbzero.debug_overlay.vplaneX[-1] ;
 wire \rbzero.debug_overlay.vplaneX[-2] ;
 wire \rbzero.debug_overlay.vplaneX[-3] ;
 wire \rbzero.debug_overlay.vplaneX[-4] ;
 wire \rbzero.debug_overlay.vplaneX[-5] ;
 wire \rbzero.debug_overlay.vplaneX[-6] ;
 wire \rbzero.debug_overlay.vplaneX[-7] ;
 wire \rbzero.debug_overlay.vplaneX[-8] ;
 wire \rbzero.debug_overlay.vplaneX[-9] ;
 wire \rbzero.debug_overlay.vplaneX[0] ;
 wire \rbzero.debug_overlay.vplaneX[10] ;
 wire \rbzero.debug_overlay.vplaneY[-1] ;
 wire \rbzero.debug_overlay.vplaneY[-2] ;
 wire \rbzero.debug_overlay.vplaneY[-3] ;
 wire \rbzero.debug_overlay.vplaneY[-4] ;
 wire \rbzero.debug_overlay.vplaneY[-5] ;
 wire \rbzero.debug_overlay.vplaneY[-6] ;
 wire \rbzero.debug_overlay.vplaneY[-7] ;
 wire \rbzero.debug_overlay.vplaneY[-8] ;
 wire \rbzero.debug_overlay.vplaneY[-9] ;
 wire \rbzero.debug_overlay.vplaneY[0] ;
 wire \rbzero.debug_overlay.vplaneY[10] ;
 wire \rbzero.floor_leak[0] ;
 wire \rbzero.floor_leak[1] ;
 wire \rbzero.floor_leak[2] ;
 wire \rbzero.floor_leak[3] ;
 wire \rbzero.floor_leak[4] ;
 wire \rbzero.floor_leak[5] ;
 wire \rbzero.hsync ;
 wire \rbzero.map_overlay.i_mapdx[0] ;
 wire \rbzero.map_overlay.i_mapdx[1] ;
 wire \rbzero.map_overlay.i_mapdx[2] ;
 wire \rbzero.map_overlay.i_mapdx[3] ;
 wire \rbzero.map_overlay.i_mapdx[4] ;
 wire \rbzero.map_overlay.i_mapdx[5] ;
 wire \rbzero.map_overlay.i_mapdy[0] ;
 wire \rbzero.map_overlay.i_mapdy[1] ;
 wire \rbzero.map_overlay.i_mapdy[2] ;
 wire \rbzero.map_overlay.i_mapdy[3] ;
 wire \rbzero.map_overlay.i_mapdy[4] ;
 wire \rbzero.map_overlay.i_mapdy[5] ;
 wire \rbzero.map_overlay.i_otherx[0] ;
 wire \rbzero.map_overlay.i_otherx[1] ;
 wire \rbzero.map_overlay.i_otherx[2] ;
 wire \rbzero.map_overlay.i_otherx[3] ;
 wire \rbzero.map_overlay.i_otherx[4] ;
 wire \rbzero.map_overlay.i_othery[0] ;
 wire \rbzero.map_overlay.i_othery[1] ;
 wire \rbzero.map_overlay.i_othery[2] ;
 wire \rbzero.map_overlay.i_othery[3] ;
 wire \rbzero.map_overlay.i_othery[4] ;
 wire \rbzero.map_rom.a6 ;
 wire \rbzero.map_rom.b6 ;
 wire \rbzero.map_rom.c6 ;
 wire \rbzero.map_rom.d6 ;
 wire \rbzero.map_rom.f1 ;
 wire \rbzero.map_rom.f2 ;
 wire \rbzero.map_rom.f3 ;
 wire \rbzero.map_rom.f4 ;
 wire \rbzero.map_rom.i_col[4] ;
 wire \rbzero.map_rom.i_row[4] ;
 wire \rbzero.mapdxw[0] ;
 wire \rbzero.mapdxw[1] ;
 wire \rbzero.mapdyw[0] ;
 wire \rbzero.mapdyw[1] ;
 wire \rbzero.pov.mosi ;
 wire \rbzero.pov.mosi_buffer[0] ;
 wire \rbzero.pov.ready ;
 wire \rbzero.pov.ready_buffer[0] ;
 wire \rbzero.pov.ready_buffer[10] ;
 wire \rbzero.pov.ready_buffer[11] ;
 wire \rbzero.pov.ready_buffer[12] ;
 wire \rbzero.pov.ready_buffer[13] ;
 wire \rbzero.pov.ready_buffer[14] ;
 wire \rbzero.pov.ready_buffer[15] ;
 wire \rbzero.pov.ready_buffer[16] ;
 wire \rbzero.pov.ready_buffer[17] ;
 wire \rbzero.pov.ready_buffer[18] ;
 wire \rbzero.pov.ready_buffer[19] ;
 wire \rbzero.pov.ready_buffer[1] ;
 wire \rbzero.pov.ready_buffer[20] ;
 wire \rbzero.pov.ready_buffer[21] ;
 wire \rbzero.pov.ready_buffer[22] ;
 wire \rbzero.pov.ready_buffer[23] ;
 wire \rbzero.pov.ready_buffer[24] ;
 wire \rbzero.pov.ready_buffer[25] ;
 wire \rbzero.pov.ready_buffer[26] ;
 wire \rbzero.pov.ready_buffer[27] ;
 wire \rbzero.pov.ready_buffer[28] ;
 wire \rbzero.pov.ready_buffer[29] ;
 wire \rbzero.pov.ready_buffer[2] ;
 wire \rbzero.pov.ready_buffer[30] ;
 wire \rbzero.pov.ready_buffer[31] ;
 wire \rbzero.pov.ready_buffer[32] ;
 wire \rbzero.pov.ready_buffer[33] ;
 wire \rbzero.pov.ready_buffer[34] ;
 wire \rbzero.pov.ready_buffer[35] ;
 wire \rbzero.pov.ready_buffer[36] ;
 wire \rbzero.pov.ready_buffer[37] ;
 wire \rbzero.pov.ready_buffer[38] ;
 wire \rbzero.pov.ready_buffer[39] ;
 wire \rbzero.pov.ready_buffer[3] ;
 wire \rbzero.pov.ready_buffer[40] ;
 wire \rbzero.pov.ready_buffer[41] ;
 wire \rbzero.pov.ready_buffer[42] ;
 wire \rbzero.pov.ready_buffer[43] ;
 wire \rbzero.pov.ready_buffer[44] ;
 wire \rbzero.pov.ready_buffer[45] ;
 wire \rbzero.pov.ready_buffer[46] ;
 wire \rbzero.pov.ready_buffer[47] ;
 wire \rbzero.pov.ready_buffer[48] ;
 wire \rbzero.pov.ready_buffer[49] ;
 wire \rbzero.pov.ready_buffer[4] ;
 wire \rbzero.pov.ready_buffer[50] ;
 wire \rbzero.pov.ready_buffer[51] ;
 wire \rbzero.pov.ready_buffer[52] ;
 wire \rbzero.pov.ready_buffer[53] ;
 wire \rbzero.pov.ready_buffer[54] ;
 wire \rbzero.pov.ready_buffer[55] ;
 wire \rbzero.pov.ready_buffer[56] ;
 wire \rbzero.pov.ready_buffer[57] ;
 wire \rbzero.pov.ready_buffer[58] ;
 wire \rbzero.pov.ready_buffer[59] ;
 wire \rbzero.pov.ready_buffer[5] ;
 wire \rbzero.pov.ready_buffer[60] ;
 wire \rbzero.pov.ready_buffer[61] ;
 wire \rbzero.pov.ready_buffer[62] ;
 wire \rbzero.pov.ready_buffer[63] ;
 wire \rbzero.pov.ready_buffer[64] ;
 wire \rbzero.pov.ready_buffer[65] ;
 wire \rbzero.pov.ready_buffer[66] ;
 wire \rbzero.pov.ready_buffer[67] ;
 wire \rbzero.pov.ready_buffer[68] ;
 wire \rbzero.pov.ready_buffer[69] ;
 wire \rbzero.pov.ready_buffer[6] ;
 wire \rbzero.pov.ready_buffer[70] ;
 wire \rbzero.pov.ready_buffer[71] ;
 wire \rbzero.pov.ready_buffer[72] ;
 wire \rbzero.pov.ready_buffer[73] ;
 wire \rbzero.pov.ready_buffer[7] ;
 wire \rbzero.pov.ready_buffer[8] ;
 wire \rbzero.pov.ready_buffer[9] ;
 wire \rbzero.pov.sclk_buffer[0] ;
 wire \rbzero.pov.sclk_buffer[1] ;
 wire \rbzero.pov.sclk_buffer[2] ;
 wire \rbzero.pov.spi_buffer[0] ;
 wire \rbzero.pov.spi_buffer[10] ;
 wire \rbzero.pov.spi_buffer[11] ;
 wire \rbzero.pov.spi_buffer[12] ;
 wire \rbzero.pov.spi_buffer[13] ;
 wire \rbzero.pov.spi_buffer[14] ;
 wire \rbzero.pov.spi_buffer[15] ;
 wire \rbzero.pov.spi_buffer[16] ;
 wire \rbzero.pov.spi_buffer[17] ;
 wire \rbzero.pov.spi_buffer[18] ;
 wire \rbzero.pov.spi_buffer[19] ;
 wire \rbzero.pov.spi_buffer[1] ;
 wire \rbzero.pov.spi_buffer[20] ;
 wire \rbzero.pov.spi_buffer[21] ;
 wire \rbzero.pov.spi_buffer[22] ;
 wire \rbzero.pov.spi_buffer[23] ;
 wire \rbzero.pov.spi_buffer[24] ;
 wire \rbzero.pov.spi_buffer[25] ;
 wire \rbzero.pov.spi_buffer[26] ;
 wire \rbzero.pov.spi_buffer[27] ;
 wire \rbzero.pov.spi_buffer[28] ;
 wire \rbzero.pov.spi_buffer[29] ;
 wire \rbzero.pov.spi_buffer[2] ;
 wire \rbzero.pov.spi_buffer[30] ;
 wire \rbzero.pov.spi_buffer[31] ;
 wire \rbzero.pov.spi_buffer[32] ;
 wire \rbzero.pov.spi_buffer[33] ;
 wire \rbzero.pov.spi_buffer[34] ;
 wire \rbzero.pov.spi_buffer[35] ;
 wire \rbzero.pov.spi_buffer[36] ;
 wire \rbzero.pov.spi_buffer[37] ;
 wire \rbzero.pov.spi_buffer[38] ;
 wire \rbzero.pov.spi_buffer[39] ;
 wire \rbzero.pov.spi_buffer[3] ;
 wire \rbzero.pov.spi_buffer[40] ;
 wire \rbzero.pov.spi_buffer[41] ;
 wire \rbzero.pov.spi_buffer[42] ;
 wire \rbzero.pov.spi_buffer[43] ;
 wire \rbzero.pov.spi_buffer[44] ;
 wire \rbzero.pov.spi_buffer[45] ;
 wire \rbzero.pov.spi_buffer[46] ;
 wire \rbzero.pov.spi_buffer[47] ;
 wire \rbzero.pov.spi_buffer[48] ;
 wire \rbzero.pov.spi_buffer[49] ;
 wire \rbzero.pov.spi_buffer[4] ;
 wire \rbzero.pov.spi_buffer[50] ;
 wire \rbzero.pov.spi_buffer[51] ;
 wire \rbzero.pov.spi_buffer[52] ;
 wire \rbzero.pov.spi_buffer[53] ;
 wire \rbzero.pov.spi_buffer[54] ;
 wire \rbzero.pov.spi_buffer[55] ;
 wire \rbzero.pov.spi_buffer[56] ;
 wire \rbzero.pov.spi_buffer[57] ;
 wire \rbzero.pov.spi_buffer[58] ;
 wire \rbzero.pov.spi_buffer[59] ;
 wire \rbzero.pov.spi_buffer[5] ;
 wire \rbzero.pov.spi_buffer[60] ;
 wire \rbzero.pov.spi_buffer[61] ;
 wire \rbzero.pov.spi_buffer[62] ;
 wire \rbzero.pov.spi_buffer[63] ;
 wire \rbzero.pov.spi_buffer[64] ;
 wire \rbzero.pov.spi_buffer[65] ;
 wire \rbzero.pov.spi_buffer[66] ;
 wire \rbzero.pov.spi_buffer[67] ;
 wire \rbzero.pov.spi_buffer[68] ;
 wire \rbzero.pov.spi_buffer[69] ;
 wire \rbzero.pov.spi_buffer[6] ;
 wire \rbzero.pov.spi_buffer[70] ;
 wire \rbzero.pov.spi_buffer[71] ;
 wire \rbzero.pov.spi_buffer[72] ;
 wire \rbzero.pov.spi_buffer[73] ;
 wire \rbzero.pov.spi_buffer[7] ;
 wire \rbzero.pov.spi_buffer[8] ;
 wire \rbzero.pov.spi_buffer[9] ;
 wire \rbzero.pov.spi_counter[0] ;
 wire \rbzero.pov.spi_counter[1] ;
 wire \rbzero.pov.spi_counter[2] ;
 wire \rbzero.pov.spi_counter[3] ;
 wire \rbzero.pov.spi_counter[4] ;
 wire \rbzero.pov.spi_counter[5] ;
 wire \rbzero.pov.spi_counter[6] ;
 wire \rbzero.pov.spi_done ;
 wire \rbzero.pov.ss_buffer[0] ;
 wire \rbzero.pov.ss_buffer[1] ;
 wire \rbzero.row_render.side ;
 wire \rbzero.row_render.size[0] ;
 wire \rbzero.row_render.size[10] ;
 wire \rbzero.row_render.size[1] ;
 wire \rbzero.row_render.size[2] ;
 wire \rbzero.row_render.size[3] ;
 wire \rbzero.row_render.size[4] ;
 wire \rbzero.row_render.size[5] ;
 wire \rbzero.row_render.size[6] ;
 wire \rbzero.row_render.size[7] ;
 wire \rbzero.row_render.size[8] ;
 wire \rbzero.row_render.size[9] ;
 wire \rbzero.row_render.texu[0] ;
 wire \rbzero.row_render.texu[1] ;
 wire \rbzero.row_render.texu[2] ;
 wire \rbzero.row_render.texu[3] ;
 wire \rbzero.row_render.texu[4] ;
 wire \rbzero.row_render.vinf ;
 wire \rbzero.row_render.wall[0] ;
 wire \rbzero.row_render.wall[1] ;
 wire \rbzero.side_hot ;
 wire \rbzero.spi_registers.got_new_floor ;
 wire \rbzero.spi_registers.got_new_leak ;
 wire \rbzero.spi_registers.got_new_mapd ;
 wire \rbzero.spi_registers.got_new_other ;
 wire \rbzero.spi_registers.got_new_sky ;
 wire \rbzero.spi_registers.got_new_texadd[0] ;
 wire \rbzero.spi_registers.got_new_texadd[1] ;
 wire \rbzero.spi_registers.got_new_texadd[2] ;
 wire \rbzero.spi_registers.got_new_texadd[3] ;
 wire \rbzero.spi_registers.got_new_vinf ;
 wire \rbzero.spi_registers.got_new_vshift ;
 wire \rbzero.spi_registers.mosi ;
 wire \rbzero.spi_registers.mosi_buffer[0] ;
 wire \rbzero.spi_registers.new_floor[0] ;
 wire \rbzero.spi_registers.new_floor[1] ;
 wire \rbzero.spi_registers.new_floor[2] ;
 wire \rbzero.spi_registers.new_floor[3] ;
 wire \rbzero.spi_registers.new_floor[4] ;
 wire \rbzero.spi_registers.new_floor[5] ;
 wire \rbzero.spi_registers.new_leak[0] ;
 wire \rbzero.spi_registers.new_leak[1] ;
 wire \rbzero.spi_registers.new_leak[2] ;
 wire \rbzero.spi_registers.new_leak[3] ;
 wire \rbzero.spi_registers.new_leak[4] ;
 wire \rbzero.spi_registers.new_leak[5] ;
 wire \rbzero.spi_registers.new_mapd[0] ;
 wire \rbzero.spi_registers.new_mapd[10] ;
 wire \rbzero.spi_registers.new_mapd[11] ;
 wire \rbzero.spi_registers.new_mapd[12] ;
 wire \rbzero.spi_registers.new_mapd[13] ;
 wire \rbzero.spi_registers.new_mapd[14] ;
 wire \rbzero.spi_registers.new_mapd[15] ;
 wire \rbzero.spi_registers.new_mapd[1] ;
 wire \rbzero.spi_registers.new_mapd[2] ;
 wire \rbzero.spi_registers.new_mapd[3] ;
 wire \rbzero.spi_registers.new_mapd[4] ;
 wire \rbzero.spi_registers.new_mapd[5] ;
 wire \rbzero.spi_registers.new_mapd[6] ;
 wire \rbzero.spi_registers.new_mapd[7] ;
 wire \rbzero.spi_registers.new_mapd[8] ;
 wire \rbzero.spi_registers.new_mapd[9] ;
 wire \rbzero.spi_registers.new_other[0] ;
 wire \rbzero.spi_registers.new_other[10] ;
 wire \rbzero.spi_registers.new_other[1] ;
 wire \rbzero.spi_registers.new_other[2] ;
 wire \rbzero.spi_registers.new_other[3] ;
 wire \rbzero.spi_registers.new_other[4] ;
 wire \rbzero.spi_registers.new_other[6] ;
 wire \rbzero.spi_registers.new_other[7] ;
 wire \rbzero.spi_registers.new_other[8] ;
 wire \rbzero.spi_registers.new_other[9] ;
 wire \rbzero.spi_registers.new_sky[0] ;
 wire \rbzero.spi_registers.new_sky[1] ;
 wire \rbzero.spi_registers.new_sky[2] ;
 wire \rbzero.spi_registers.new_sky[3] ;
 wire \rbzero.spi_registers.new_sky[4] ;
 wire \rbzero.spi_registers.new_sky[5] ;
 wire \rbzero.spi_registers.new_texadd[0][0] ;
 wire \rbzero.spi_registers.new_texadd[0][10] ;
 wire \rbzero.spi_registers.new_texadd[0][11] ;
 wire \rbzero.spi_registers.new_texadd[0][12] ;
 wire \rbzero.spi_registers.new_texadd[0][13] ;
 wire \rbzero.spi_registers.new_texadd[0][14] ;
 wire \rbzero.spi_registers.new_texadd[0][15] ;
 wire \rbzero.spi_registers.new_texadd[0][16] ;
 wire \rbzero.spi_registers.new_texadd[0][17] ;
 wire \rbzero.spi_registers.new_texadd[0][18] ;
 wire \rbzero.spi_registers.new_texadd[0][19] ;
 wire \rbzero.spi_registers.new_texadd[0][1] ;
 wire \rbzero.spi_registers.new_texadd[0][20] ;
 wire \rbzero.spi_registers.new_texadd[0][21] ;
 wire \rbzero.spi_registers.new_texadd[0][22] ;
 wire \rbzero.spi_registers.new_texadd[0][23] ;
 wire \rbzero.spi_registers.new_texadd[0][2] ;
 wire \rbzero.spi_registers.new_texadd[0][3] ;
 wire \rbzero.spi_registers.new_texadd[0][4] ;
 wire \rbzero.spi_registers.new_texadd[0][5] ;
 wire \rbzero.spi_registers.new_texadd[0][6] ;
 wire \rbzero.spi_registers.new_texadd[0][7] ;
 wire \rbzero.spi_registers.new_texadd[0][8] ;
 wire \rbzero.spi_registers.new_texadd[0][9] ;
 wire \rbzero.spi_registers.new_texadd[1][0] ;
 wire \rbzero.spi_registers.new_texadd[1][10] ;
 wire \rbzero.spi_registers.new_texadd[1][11] ;
 wire \rbzero.spi_registers.new_texadd[1][12] ;
 wire \rbzero.spi_registers.new_texadd[1][13] ;
 wire \rbzero.spi_registers.new_texadd[1][14] ;
 wire \rbzero.spi_registers.new_texadd[1][15] ;
 wire \rbzero.spi_registers.new_texadd[1][16] ;
 wire \rbzero.spi_registers.new_texadd[1][17] ;
 wire \rbzero.spi_registers.new_texadd[1][18] ;
 wire \rbzero.spi_registers.new_texadd[1][19] ;
 wire \rbzero.spi_registers.new_texadd[1][1] ;
 wire \rbzero.spi_registers.new_texadd[1][20] ;
 wire \rbzero.spi_registers.new_texadd[1][21] ;
 wire \rbzero.spi_registers.new_texadd[1][22] ;
 wire \rbzero.spi_registers.new_texadd[1][23] ;
 wire \rbzero.spi_registers.new_texadd[1][2] ;
 wire \rbzero.spi_registers.new_texadd[1][3] ;
 wire \rbzero.spi_registers.new_texadd[1][4] ;
 wire \rbzero.spi_registers.new_texadd[1][5] ;
 wire \rbzero.spi_registers.new_texadd[1][6] ;
 wire \rbzero.spi_registers.new_texadd[1][7] ;
 wire \rbzero.spi_registers.new_texadd[1][8] ;
 wire \rbzero.spi_registers.new_texadd[1][9] ;
 wire \rbzero.spi_registers.new_texadd[2][0] ;
 wire \rbzero.spi_registers.new_texadd[2][10] ;
 wire \rbzero.spi_registers.new_texadd[2][11] ;
 wire \rbzero.spi_registers.new_texadd[2][12] ;
 wire \rbzero.spi_registers.new_texadd[2][13] ;
 wire \rbzero.spi_registers.new_texadd[2][14] ;
 wire \rbzero.spi_registers.new_texadd[2][15] ;
 wire \rbzero.spi_registers.new_texadd[2][16] ;
 wire \rbzero.spi_registers.new_texadd[2][17] ;
 wire \rbzero.spi_registers.new_texadd[2][18] ;
 wire \rbzero.spi_registers.new_texadd[2][19] ;
 wire \rbzero.spi_registers.new_texadd[2][1] ;
 wire \rbzero.spi_registers.new_texadd[2][20] ;
 wire \rbzero.spi_registers.new_texadd[2][21] ;
 wire \rbzero.spi_registers.new_texadd[2][22] ;
 wire \rbzero.spi_registers.new_texadd[2][23] ;
 wire \rbzero.spi_registers.new_texadd[2][2] ;
 wire \rbzero.spi_registers.new_texadd[2][3] ;
 wire \rbzero.spi_registers.new_texadd[2][4] ;
 wire \rbzero.spi_registers.new_texadd[2][5] ;
 wire \rbzero.spi_registers.new_texadd[2][6] ;
 wire \rbzero.spi_registers.new_texadd[2][7] ;
 wire \rbzero.spi_registers.new_texadd[2][8] ;
 wire \rbzero.spi_registers.new_texadd[2][9] ;
 wire \rbzero.spi_registers.new_texadd[3][0] ;
 wire \rbzero.spi_registers.new_texadd[3][10] ;
 wire \rbzero.spi_registers.new_texadd[3][11] ;
 wire \rbzero.spi_registers.new_texadd[3][12] ;
 wire \rbzero.spi_registers.new_texadd[3][13] ;
 wire \rbzero.spi_registers.new_texadd[3][14] ;
 wire \rbzero.spi_registers.new_texadd[3][15] ;
 wire \rbzero.spi_registers.new_texadd[3][16] ;
 wire \rbzero.spi_registers.new_texadd[3][17] ;
 wire \rbzero.spi_registers.new_texadd[3][18] ;
 wire \rbzero.spi_registers.new_texadd[3][19] ;
 wire \rbzero.spi_registers.new_texadd[3][1] ;
 wire \rbzero.spi_registers.new_texadd[3][20] ;
 wire \rbzero.spi_registers.new_texadd[3][21] ;
 wire \rbzero.spi_registers.new_texadd[3][22] ;
 wire \rbzero.spi_registers.new_texadd[3][23] ;
 wire \rbzero.spi_registers.new_texadd[3][2] ;
 wire \rbzero.spi_registers.new_texadd[3][3] ;
 wire \rbzero.spi_registers.new_texadd[3][4] ;
 wire \rbzero.spi_registers.new_texadd[3][5] ;
 wire \rbzero.spi_registers.new_texadd[3][6] ;
 wire \rbzero.spi_registers.new_texadd[3][7] ;
 wire \rbzero.spi_registers.new_texadd[3][8] ;
 wire \rbzero.spi_registers.new_texadd[3][9] ;
 wire \rbzero.spi_registers.new_vinf ;
 wire \rbzero.spi_registers.new_vshift[0] ;
 wire \rbzero.spi_registers.new_vshift[1] ;
 wire \rbzero.spi_registers.new_vshift[2] ;
 wire \rbzero.spi_registers.new_vshift[3] ;
 wire \rbzero.spi_registers.new_vshift[4] ;
 wire \rbzero.spi_registers.new_vshift[5] ;
 wire \rbzero.spi_registers.sclk_buffer[0] ;
 wire \rbzero.spi_registers.sclk_buffer[1] ;
 wire \rbzero.spi_registers.sclk_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[0] ;
 wire \rbzero.spi_registers.spi_buffer[10] ;
 wire \rbzero.spi_registers.spi_buffer[11] ;
 wire \rbzero.spi_registers.spi_buffer[12] ;
 wire \rbzero.spi_registers.spi_buffer[13] ;
 wire \rbzero.spi_registers.spi_buffer[14] ;
 wire \rbzero.spi_registers.spi_buffer[15] ;
 wire \rbzero.spi_registers.spi_buffer[16] ;
 wire \rbzero.spi_registers.spi_buffer[17] ;
 wire \rbzero.spi_registers.spi_buffer[18] ;
 wire \rbzero.spi_registers.spi_buffer[19] ;
 wire \rbzero.spi_registers.spi_buffer[1] ;
 wire \rbzero.spi_registers.spi_buffer[20] ;
 wire \rbzero.spi_registers.spi_buffer[21] ;
 wire \rbzero.spi_registers.spi_buffer[22] ;
 wire \rbzero.spi_registers.spi_buffer[23] ;
 wire \rbzero.spi_registers.spi_buffer[2] ;
 wire \rbzero.spi_registers.spi_buffer[3] ;
 wire \rbzero.spi_registers.spi_buffer[4] ;
 wire \rbzero.spi_registers.spi_buffer[5] ;
 wire \rbzero.spi_registers.spi_buffer[6] ;
 wire \rbzero.spi_registers.spi_buffer[7] ;
 wire \rbzero.spi_registers.spi_buffer[8] ;
 wire \rbzero.spi_registers.spi_buffer[9] ;
 wire \rbzero.spi_registers.spi_cmd[0] ;
 wire \rbzero.spi_registers.spi_cmd[1] ;
 wire \rbzero.spi_registers.spi_cmd[2] ;
 wire \rbzero.spi_registers.spi_cmd[3] ;
 wire \rbzero.spi_registers.spi_counter[0] ;
 wire \rbzero.spi_registers.spi_counter[1] ;
 wire \rbzero.spi_registers.spi_counter[2] ;
 wire \rbzero.spi_registers.spi_counter[3] ;
 wire \rbzero.spi_registers.spi_counter[4] ;
 wire \rbzero.spi_registers.spi_counter[5] ;
 wire \rbzero.spi_registers.spi_counter[6] ;
 wire \rbzero.spi_registers.spi_done ;
 wire \rbzero.spi_registers.ss_buffer[0] ;
 wire \rbzero.spi_registers.ss_buffer[1] ;
 wire \rbzero.spi_registers.texadd0[0] ;
 wire \rbzero.spi_registers.texadd0[10] ;
 wire \rbzero.spi_registers.texadd0[11] ;
 wire \rbzero.spi_registers.texadd0[12] ;
 wire \rbzero.spi_registers.texadd0[13] ;
 wire \rbzero.spi_registers.texadd0[14] ;
 wire \rbzero.spi_registers.texadd0[15] ;
 wire \rbzero.spi_registers.texadd0[16] ;
 wire \rbzero.spi_registers.texadd0[17] ;
 wire \rbzero.spi_registers.texadd0[18] ;
 wire \rbzero.spi_registers.texadd0[19] ;
 wire \rbzero.spi_registers.texadd0[1] ;
 wire \rbzero.spi_registers.texadd0[20] ;
 wire \rbzero.spi_registers.texadd0[21] ;
 wire \rbzero.spi_registers.texadd0[22] ;
 wire \rbzero.spi_registers.texadd0[23] ;
 wire \rbzero.spi_registers.texadd0[2] ;
 wire \rbzero.spi_registers.texadd0[3] ;
 wire \rbzero.spi_registers.texadd0[4] ;
 wire \rbzero.spi_registers.texadd0[5] ;
 wire \rbzero.spi_registers.texadd0[6] ;
 wire \rbzero.spi_registers.texadd0[7] ;
 wire \rbzero.spi_registers.texadd0[8] ;
 wire \rbzero.spi_registers.texadd0[9] ;
 wire \rbzero.spi_registers.texadd1[0] ;
 wire \rbzero.spi_registers.texadd1[10] ;
 wire \rbzero.spi_registers.texadd1[11] ;
 wire \rbzero.spi_registers.texadd1[12] ;
 wire \rbzero.spi_registers.texadd1[13] ;
 wire \rbzero.spi_registers.texadd1[14] ;
 wire \rbzero.spi_registers.texadd1[15] ;
 wire \rbzero.spi_registers.texadd1[16] ;
 wire \rbzero.spi_registers.texadd1[17] ;
 wire \rbzero.spi_registers.texadd1[18] ;
 wire \rbzero.spi_registers.texadd1[19] ;
 wire \rbzero.spi_registers.texadd1[1] ;
 wire \rbzero.spi_registers.texadd1[20] ;
 wire \rbzero.spi_registers.texadd1[21] ;
 wire \rbzero.spi_registers.texadd1[22] ;
 wire \rbzero.spi_registers.texadd1[23] ;
 wire \rbzero.spi_registers.texadd1[2] ;
 wire \rbzero.spi_registers.texadd1[3] ;
 wire \rbzero.spi_registers.texadd1[4] ;
 wire \rbzero.spi_registers.texadd1[5] ;
 wire \rbzero.spi_registers.texadd1[6] ;
 wire \rbzero.spi_registers.texadd1[7] ;
 wire \rbzero.spi_registers.texadd1[8] ;
 wire \rbzero.spi_registers.texadd1[9] ;
 wire \rbzero.spi_registers.texadd2[0] ;
 wire \rbzero.spi_registers.texadd2[10] ;
 wire \rbzero.spi_registers.texadd2[11] ;
 wire \rbzero.spi_registers.texadd2[12] ;
 wire \rbzero.spi_registers.texadd2[13] ;
 wire \rbzero.spi_registers.texadd2[14] ;
 wire \rbzero.spi_registers.texadd2[15] ;
 wire \rbzero.spi_registers.texadd2[16] ;
 wire \rbzero.spi_registers.texadd2[17] ;
 wire \rbzero.spi_registers.texadd2[18] ;
 wire \rbzero.spi_registers.texadd2[19] ;
 wire \rbzero.spi_registers.texadd2[1] ;
 wire \rbzero.spi_registers.texadd2[20] ;
 wire \rbzero.spi_registers.texadd2[21] ;
 wire \rbzero.spi_registers.texadd2[22] ;
 wire \rbzero.spi_registers.texadd2[23] ;
 wire \rbzero.spi_registers.texadd2[2] ;
 wire \rbzero.spi_registers.texadd2[3] ;
 wire \rbzero.spi_registers.texadd2[4] ;
 wire \rbzero.spi_registers.texadd2[5] ;
 wire \rbzero.spi_registers.texadd2[6] ;
 wire \rbzero.spi_registers.texadd2[7] ;
 wire \rbzero.spi_registers.texadd2[8] ;
 wire \rbzero.spi_registers.texadd2[9] ;
 wire \rbzero.spi_registers.texadd3[0] ;
 wire \rbzero.spi_registers.texadd3[10] ;
 wire \rbzero.spi_registers.texadd3[11] ;
 wire \rbzero.spi_registers.texadd3[12] ;
 wire \rbzero.spi_registers.texadd3[13] ;
 wire \rbzero.spi_registers.texadd3[14] ;
 wire \rbzero.spi_registers.texadd3[15] ;
 wire \rbzero.spi_registers.texadd3[16] ;
 wire \rbzero.spi_registers.texadd3[17] ;
 wire \rbzero.spi_registers.texadd3[18] ;
 wire \rbzero.spi_registers.texadd3[19] ;
 wire \rbzero.spi_registers.texadd3[1] ;
 wire \rbzero.spi_registers.texadd3[20] ;
 wire \rbzero.spi_registers.texadd3[21] ;
 wire \rbzero.spi_registers.texadd3[22] ;
 wire \rbzero.spi_registers.texadd3[23] ;
 wire \rbzero.spi_registers.texadd3[2] ;
 wire \rbzero.spi_registers.texadd3[3] ;
 wire \rbzero.spi_registers.texadd3[4] ;
 wire \rbzero.spi_registers.texadd3[5] ;
 wire \rbzero.spi_registers.texadd3[6] ;
 wire \rbzero.spi_registers.texadd3[7] ;
 wire \rbzero.spi_registers.texadd3[8] ;
 wire \rbzero.spi_registers.texadd3[9] ;
 wire \rbzero.spi_registers.vshift[0] ;
 wire \rbzero.spi_registers.vshift[1] ;
 wire \rbzero.spi_registers.vshift[2] ;
 wire \rbzero.spi_registers.vshift[3] ;
 wire \rbzero.spi_registers.vshift[4] ;
 wire \rbzero.spi_registers.vshift[5] ;
 wire \rbzero.texV[-10] ;
 wire \rbzero.texV[-11] ;
 wire \rbzero.texV[-1] ;
 wire \rbzero.texV[-2] ;
 wire \rbzero.texV[-3] ;
 wire \rbzero.texV[-4] ;
 wire \rbzero.texV[-5] ;
 wire \rbzero.texV[-6] ;
 wire \rbzero.texV[-7] ;
 wire \rbzero.texV[-8] ;
 wire \rbzero.texV[-9] ;
 wire \rbzero.texV[0] ;
 wire \rbzero.texV[10] ;
 wire \rbzero.texV[1] ;
 wire \rbzero.texV[2] ;
 wire \rbzero.texV[3] ;
 wire \rbzero.texV[4] ;
 wire \rbzero.texV[5] ;
 wire \rbzero.texV[6] ;
 wire \rbzero.texV[7] ;
 wire \rbzero.texV[8] ;
 wire \rbzero.texV[9] ;
 wire \rbzero.tex_b0[0] ;
 wire \rbzero.tex_b0[10] ;
 wire \rbzero.tex_b0[11] ;
 wire \rbzero.tex_b0[12] ;
 wire \rbzero.tex_b0[13] ;
 wire \rbzero.tex_b0[14] ;
 wire \rbzero.tex_b0[15] ;
 wire \rbzero.tex_b0[16] ;
 wire \rbzero.tex_b0[17] ;
 wire \rbzero.tex_b0[18] ;
 wire \rbzero.tex_b0[19] ;
 wire \rbzero.tex_b0[1] ;
 wire \rbzero.tex_b0[20] ;
 wire \rbzero.tex_b0[21] ;
 wire \rbzero.tex_b0[22] ;
 wire \rbzero.tex_b0[23] ;
 wire \rbzero.tex_b0[24] ;
 wire \rbzero.tex_b0[25] ;
 wire \rbzero.tex_b0[26] ;
 wire \rbzero.tex_b0[27] ;
 wire \rbzero.tex_b0[28] ;
 wire \rbzero.tex_b0[29] ;
 wire \rbzero.tex_b0[2] ;
 wire \rbzero.tex_b0[30] ;
 wire \rbzero.tex_b0[31] ;
 wire \rbzero.tex_b0[32] ;
 wire \rbzero.tex_b0[33] ;
 wire \rbzero.tex_b0[34] ;
 wire \rbzero.tex_b0[35] ;
 wire \rbzero.tex_b0[36] ;
 wire \rbzero.tex_b0[37] ;
 wire \rbzero.tex_b0[38] ;
 wire \rbzero.tex_b0[39] ;
 wire \rbzero.tex_b0[3] ;
 wire \rbzero.tex_b0[40] ;
 wire \rbzero.tex_b0[41] ;
 wire \rbzero.tex_b0[42] ;
 wire \rbzero.tex_b0[43] ;
 wire \rbzero.tex_b0[44] ;
 wire \rbzero.tex_b0[45] ;
 wire \rbzero.tex_b0[46] ;
 wire \rbzero.tex_b0[47] ;
 wire \rbzero.tex_b0[48] ;
 wire \rbzero.tex_b0[49] ;
 wire \rbzero.tex_b0[4] ;
 wire \rbzero.tex_b0[50] ;
 wire \rbzero.tex_b0[51] ;
 wire \rbzero.tex_b0[52] ;
 wire \rbzero.tex_b0[53] ;
 wire \rbzero.tex_b0[54] ;
 wire \rbzero.tex_b0[55] ;
 wire \rbzero.tex_b0[56] ;
 wire \rbzero.tex_b0[57] ;
 wire \rbzero.tex_b0[58] ;
 wire \rbzero.tex_b0[59] ;
 wire \rbzero.tex_b0[5] ;
 wire \rbzero.tex_b0[60] ;
 wire \rbzero.tex_b0[61] ;
 wire \rbzero.tex_b0[62] ;
 wire \rbzero.tex_b0[63] ;
 wire \rbzero.tex_b0[6] ;
 wire \rbzero.tex_b0[7] ;
 wire \rbzero.tex_b0[8] ;
 wire \rbzero.tex_b0[9] ;
 wire \rbzero.tex_b1[0] ;
 wire \rbzero.tex_b1[10] ;
 wire \rbzero.tex_b1[11] ;
 wire \rbzero.tex_b1[12] ;
 wire \rbzero.tex_b1[13] ;
 wire \rbzero.tex_b1[14] ;
 wire \rbzero.tex_b1[15] ;
 wire \rbzero.tex_b1[16] ;
 wire \rbzero.tex_b1[17] ;
 wire \rbzero.tex_b1[18] ;
 wire \rbzero.tex_b1[19] ;
 wire \rbzero.tex_b1[1] ;
 wire \rbzero.tex_b1[20] ;
 wire \rbzero.tex_b1[21] ;
 wire \rbzero.tex_b1[22] ;
 wire \rbzero.tex_b1[23] ;
 wire \rbzero.tex_b1[24] ;
 wire \rbzero.tex_b1[25] ;
 wire \rbzero.tex_b1[26] ;
 wire \rbzero.tex_b1[27] ;
 wire \rbzero.tex_b1[28] ;
 wire \rbzero.tex_b1[29] ;
 wire \rbzero.tex_b1[2] ;
 wire \rbzero.tex_b1[30] ;
 wire \rbzero.tex_b1[31] ;
 wire \rbzero.tex_b1[32] ;
 wire \rbzero.tex_b1[33] ;
 wire \rbzero.tex_b1[34] ;
 wire \rbzero.tex_b1[35] ;
 wire \rbzero.tex_b1[36] ;
 wire \rbzero.tex_b1[37] ;
 wire \rbzero.tex_b1[38] ;
 wire \rbzero.tex_b1[39] ;
 wire \rbzero.tex_b1[3] ;
 wire \rbzero.tex_b1[40] ;
 wire \rbzero.tex_b1[41] ;
 wire \rbzero.tex_b1[42] ;
 wire \rbzero.tex_b1[43] ;
 wire \rbzero.tex_b1[44] ;
 wire \rbzero.tex_b1[45] ;
 wire \rbzero.tex_b1[46] ;
 wire \rbzero.tex_b1[47] ;
 wire \rbzero.tex_b1[48] ;
 wire \rbzero.tex_b1[49] ;
 wire \rbzero.tex_b1[4] ;
 wire \rbzero.tex_b1[50] ;
 wire \rbzero.tex_b1[51] ;
 wire \rbzero.tex_b1[52] ;
 wire \rbzero.tex_b1[53] ;
 wire \rbzero.tex_b1[54] ;
 wire \rbzero.tex_b1[55] ;
 wire \rbzero.tex_b1[56] ;
 wire \rbzero.tex_b1[57] ;
 wire \rbzero.tex_b1[58] ;
 wire \rbzero.tex_b1[59] ;
 wire \rbzero.tex_b1[5] ;
 wire \rbzero.tex_b1[60] ;
 wire \rbzero.tex_b1[61] ;
 wire \rbzero.tex_b1[62] ;
 wire \rbzero.tex_b1[63] ;
 wire \rbzero.tex_b1[6] ;
 wire \rbzero.tex_b1[7] ;
 wire \rbzero.tex_b1[8] ;
 wire \rbzero.tex_b1[9] ;
 wire \rbzero.tex_g0[0] ;
 wire \rbzero.tex_g0[10] ;
 wire \rbzero.tex_g0[11] ;
 wire \rbzero.tex_g0[12] ;
 wire \rbzero.tex_g0[13] ;
 wire \rbzero.tex_g0[14] ;
 wire \rbzero.tex_g0[15] ;
 wire \rbzero.tex_g0[16] ;
 wire \rbzero.tex_g0[17] ;
 wire \rbzero.tex_g0[18] ;
 wire \rbzero.tex_g0[19] ;
 wire \rbzero.tex_g0[1] ;
 wire \rbzero.tex_g0[20] ;
 wire \rbzero.tex_g0[21] ;
 wire \rbzero.tex_g0[22] ;
 wire \rbzero.tex_g0[23] ;
 wire \rbzero.tex_g0[24] ;
 wire \rbzero.tex_g0[25] ;
 wire \rbzero.tex_g0[26] ;
 wire \rbzero.tex_g0[27] ;
 wire \rbzero.tex_g0[28] ;
 wire \rbzero.tex_g0[29] ;
 wire \rbzero.tex_g0[2] ;
 wire \rbzero.tex_g0[30] ;
 wire \rbzero.tex_g0[31] ;
 wire \rbzero.tex_g0[32] ;
 wire \rbzero.tex_g0[33] ;
 wire \rbzero.tex_g0[34] ;
 wire \rbzero.tex_g0[35] ;
 wire \rbzero.tex_g0[36] ;
 wire \rbzero.tex_g0[37] ;
 wire \rbzero.tex_g0[38] ;
 wire \rbzero.tex_g0[39] ;
 wire \rbzero.tex_g0[3] ;
 wire \rbzero.tex_g0[40] ;
 wire \rbzero.tex_g0[41] ;
 wire \rbzero.tex_g0[42] ;
 wire \rbzero.tex_g0[43] ;
 wire \rbzero.tex_g0[44] ;
 wire \rbzero.tex_g0[45] ;
 wire \rbzero.tex_g0[46] ;
 wire \rbzero.tex_g0[47] ;
 wire \rbzero.tex_g0[48] ;
 wire \rbzero.tex_g0[49] ;
 wire \rbzero.tex_g0[4] ;
 wire \rbzero.tex_g0[50] ;
 wire \rbzero.tex_g0[51] ;
 wire \rbzero.tex_g0[52] ;
 wire \rbzero.tex_g0[53] ;
 wire \rbzero.tex_g0[54] ;
 wire \rbzero.tex_g0[55] ;
 wire \rbzero.tex_g0[56] ;
 wire \rbzero.tex_g0[57] ;
 wire \rbzero.tex_g0[58] ;
 wire \rbzero.tex_g0[59] ;
 wire \rbzero.tex_g0[5] ;
 wire \rbzero.tex_g0[60] ;
 wire \rbzero.tex_g0[61] ;
 wire \rbzero.tex_g0[62] ;
 wire \rbzero.tex_g0[63] ;
 wire \rbzero.tex_g0[6] ;
 wire \rbzero.tex_g0[7] ;
 wire \rbzero.tex_g0[8] ;
 wire \rbzero.tex_g0[9] ;
 wire \rbzero.tex_g1[0] ;
 wire \rbzero.tex_g1[10] ;
 wire \rbzero.tex_g1[11] ;
 wire \rbzero.tex_g1[12] ;
 wire \rbzero.tex_g1[13] ;
 wire \rbzero.tex_g1[14] ;
 wire \rbzero.tex_g1[15] ;
 wire \rbzero.tex_g1[16] ;
 wire \rbzero.tex_g1[17] ;
 wire \rbzero.tex_g1[18] ;
 wire \rbzero.tex_g1[19] ;
 wire \rbzero.tex_g1[1] ;
 wire \rbzero.tex_g1[20] ;
 wire \rbzero.tex_g1[21] ;
 wire \rbzero.tex_g1[22] ;
 wire \rbzero.tex_g1[23] ;
 wire \rbzero.tex_g1[24] ;
 wire \rbzero.tex_g1[25] ;
 wire \rbzero.tex_g1[26] ;
 wire \rbzero.tex_g1[27] ;
 wire \rbzero.tex_g1[28] ;
 wire \rbzero.tex_g1[29] ;
 wire \rbzero.tex_g1[2] ;
 wire \rbzero.tex_g1[30] ;
 wire \rbzero.tex_g1[31] ;
 wire \rbzero.tex_g1[32] ;
 wire \rbzero.tex_g1[33] ;
 wire \rbzero.tex_g1[34] ;
 wire \rbzero.tex_g1[35] ;
 wire \rbzero.tex_g1[36] ;
 wire \rbzero.tex_g1[37] ;
 wire \rbzero.tex_g1[38] ;
 wire \rbzero.tex_g1[39] ;
 wire \rbzero.tex_g1[3] ;
 wire \rbzero.tex_g1[40] ;
 wire \rbzero.tex_g1[41] ;
 wire \rbzero.tex_g1[42] ;
 wire \rbzero.tex_g1[43] ;
 wire \rbzero.tex_g1[44] ;
 wire \rbzero.tex_g1[45] ;
 wire \rbzero.tex_g1[46] ;
 wire \rbzero.tex_g1[47] ;
 wire \rbzero.tex_g1[48] ;
 wire \rbzero.tex_g1[49] ;
 wire \rbzero.tex_g1[4] ;
 wire \rbzero.tex_g1[50] ;
 wire \rbzero.tex_g1[51] ;
 wire \rbzero.tex_g1[52] ;
 wire \rbzero.tex_g1[53] ;
 wire \rbzero.tex_g1[54] ;
 wire \rbzero.tex_g1[55] ;
 wire \rbzero.tex_g1[56] ;
 wire \rbzero.tex_g1[57] ;
 wire \rbzero.tex_g1[58] ;
 wire \rbzero.tex_g1[59] ;
 wire \rbzero.tex_g1[5] ;
 wire \rbzero.tex_g1[60] ;
 wire \rbzero.tex_g1[61] ;
 wire \rbzero.tex_g1[62] ;
 wire \rbzero.tex_g1[63] ;
 wire \rbzero.tex_g1[6] ;
 wire \rbzero.tex_g1[7] ;
 wire \rbzero.tex_g1[8] ;
 wire \rbzero.tex_g1[9] ;
 wire \rbzero.tex_r0[0] ;
 wire \rbzero.tex_r0[10] ;
 wire \rbzero.tex_r0[11] ;
 wire \rbzero.tex_r0[12] ;
 wire \rbzero.tex_r0[13] ;
 wire \rbzero.tex_r0[14] ;
 wire \rbzero.tex_r0[15] ;
 wire \rbzero.tex_r0[16] ;
 wire \rbzero.tex_r0[17] ;
 wire \rbzero.tex_r0[18] ;
 wire \rbzero.tex_r0[19] ;
 wire \rbzero.tex_r0[1] ;
 wire \rbzero.tex_r0[20] ;
 wire \rbzero.tex_r0[21] ;
 wire \rbzero.tex_r0[22] ;
 wire \rbzero.tex_r0[23] ;
 wire \rbzero.tex_r0[24] ;
 wire \rbzero.tex_r0[25] ;
 wire \rbzero.tex_r0[26] ;
 wire \rbzero.tex_r0[27] ;
 wire \rbzero.tex_r0[28] ;
 wire \rbzero.tex_r0[29] ;
 wire \rbzero.tex_r0[2] ;
 wire \rbzero.tex_r0[30] ;
 wire \rbzero.tex_r0[31] ;
 wire \rbzero.tex_r0[32] ;
 wire \rbzero.tex_r0[33] ;
 wire \rbzero.tex_r0[34] ;
 wire \rbzero.tex_r0[35] ;
 wire \rbzero.tex_r0[36] ;
 wire \rbzero.tex_r0[37] ;
 wire \rbzero.tex_r0[38] ;
 wire \rbzero.tex_r0[39] ;
 wire \rbzero.tex_r0[3] ;
 wire \rbzero.tex_r0[40] ;
 wire \rbzero.tex_r0[41] ;
 wire \rbzero.tex_r0[42] ;
 wire \rbzero.tex_r0[43] ;
 wire \rbzero.tex_r0[44] ;
 wire \rbzero.tex_r0[45] ;
 wire \rbzero.tex_r0[46] ;
 wire \rbzero.tex_r0[47] ;
 wire \rbzero.tex_r0[48] ;
 wire \rbzero.tex_r0[49] ;
 wire \rbzero.tex_r0[4] ;
 wire \rbzero.tex_r0[50] ;
 wire \rbzero.tex_r0[51] ;
 wire \rbzero.tex_r0[52] ;
 wire \rbzero.tex_r0[53] ;
 wire \rbzero.tex_r0[54] ;
 wire \rbzero.tex_r0[55] ;
 wire \rbzero.tex_r0[56] ;
 wire \rbzero.tex_r0[57] ;
 wire \rbzero.tex_r0[58] ;
 wire \rbzero.tex_r0[59] ;
 wire \rbzero.tex_r0[5] ;
 wire \rbzero.tex_r0[60] ;
 wire \rbzero.tex_r0[61] ;
 wire \rbzero.tex_r0[62] ;
 wire \rbzero.tex_r0[63] ;
 wire \rbzero.tex_r0[6] ;
 wire \rbzero.tex_r0[7] ;
 wire \rbzero.tex_r0[8] ;
 wire \rbzero.tex_r0[9] ;
 wire \rbzero.tex_r1[0] ;
 wire \rbzero.tex_r1[10] ;
 wire \rbzero.tex_r1[11] ;
 wire \rbzero.tex_r1[12] ;
 wire \rbzero.tex_r1[13] ;
 wire \rbzero.tex_r1[14] ;
 wire \rbzero.tex_r1[15] ;
 wire \rbzero.tex_r1[16] ;
 wire \rbzero.tex_r1[17] ;
 wire \rbzero.tex_r1[18] ;
 wire \rbzero.tex_r1[19] ;
 wire \rbzero.tex_r1[1] ;
 wire \rbzero.tex_r1[20] ;
 wire \rbzero.tex_r1[21] ;
 wire \rbzero.tex_r1[22] ;
 wire \rbzero.tex_r1[23] ;
 wire \rbzero.tex_r1[24] ;
 wire \rbzero.tex_r1[25] ;
 wire \rbzero.tex_r1[26] ;
 wire \rbzero.tex_r1[27] ;
 wire \rbzero.tex_r1[28] ;
 wire \rbzero.tex_r1[29] ;
 wire \rbzero.tex_r1[2] ;
 wire \rbzero.tex_r1[30] ;
 wire \rbzero.tex_r1[31] ;
 wire \rbzero.tex_r1[32] ;
 wire \rbzero.tex_r1[33] ;
 wire \rbzero.tex_r1[34] ;
 wire \rbzero.tex_r1[35] ;
 wire \rbzero.tex_r1[36] ;
 wire \rbzero.tex_r1[37] ;
 wire \rbzero.tex_r1[38] ;
 wire \rbzero.tex_r1[39] ;
 wire \rbzero.tex_r1[3] ;
 wire \rbzero.tex_r1[40] ;
 wire \rbzero.tex_r1[41] ;
 wire \rbzero.tex_r1[42] ;
 wire \rbzero.tex_r1[43] ;
 wire \rbzero.tex_r1[44] ;
 wire \rbzero.tex_r1[45] ;
 wire \rbzero.tex_r1[46] ;
 wire \rbzero.tex_r1[47] ;
 wire \rbzero.tex_r1[48] ;
 wire \rbzero.tex_r1[49] ;
 wire \rbzero.tex_r1[4] ;
 wire \rbzero.tex_r1[50] ;
 wire \rbzero.tex_r1[51] ;
 wire \rbzero.tex_r1[52] ;
 wire \rbzero.tex_r1[53] ;
 wire \rbzero.tex_r1[54] ;
 wire \rbzero.tex_r1[55] ;
 wire \rbzero.tex_r1[56] ;
 wire \rbzero.tex_r1[57] ;
 wire \rbzero.tex_r1[58] ;
 wire \rbzero.tex_r1[59] ;
 wire \rbzero.tex_r1[5] ;
 wire \rbzero.tex_r1[60] ;
 wire \rbzero.tex_r1[61] ;
 wire \rbzero.tex_r1[62] ;
 wire \rbzero.tex_r1[63] ;
 wire \rbzero.tex_r1[6] ;
 wire \rbzero.tex_r1[7] ;
 wire \rbzero.tex_r1[8] ;
 wire \rbzero.tex_r1[9] ;
 wire \rbzero.texu_hot[0] ;
 wire \rbzero.texu_hot[1] ;
 wire \rbzero.texu_hot[2] ;
 wire \rbzero.texu_hot[3] ;
 wire \rbzero.texu_hot[4] ;
 wire \rbzero.texu_hot[5] ;
 wire \rbzero.trace_state[0] ;
 wire \rbzero.trace_state[1] ;
 wire \rbzero.trace_state[2] ;
 wire \rbzero.trace_state[3] ;
 wire \rbzero.traced_texVinit[0] ;
 wire \rbzero.traced_texVinit[10] ;
 wire \rbzero.traced_texVinit[1] ;
 wire \rbzero.traced_texVinit[2] ;
 wire \rbzero.traced_texVinit[3] ;
 wire \rbzero.traced_texVinit[4] ;
 wire \rbzero.traced_texVinit[5] ;
 wire \rbzero.traced_texVinit[6] ;
 wire \rbzero.traced_texVinit[7] ;
 wire \rbzero.traced_texVinit[8] ;
 wire \rbzero.traced_texVinit[9] ;
 wire \rbzero.traced_texa[-10] ;
 wire \rbzero.traced_texa[-11] ;
 wire \rbzero.traced_texa[-1] ;
 wire \rbzero.traced_texa[-2] ;
 wire \rbzero.traced_texa[-3] ;
 wire \rbzero.traced_texa[-4] ;
 wire \rbzero.traced_texa[-5] ;
 wire \rbzero.traced_texa[-6] ;
 wire \rbzero.traced_texa[-7] ;
 wire \rbzero.traced_texa[-8] ;
 wire \rbzero.traced_texa[-9] ;
 wire \rbzero.traced_texa[0] ;
 wire \rbzero.traced_texa[10] ;
 wire \rbzero.traced_texa[1] ;
 wire \rbzero.traced_texa[2] ;
 wire \rbzero.traced_texa[3] ;
 wire \rbzero.traced_texa[4] ;
 wire \rbzero.traced_texa[5] ;
 wire \rbzero.traced_texa[6] ;
 wire \rbzero.traced_texa[7] ;
 wire \rbzero.traced_texa[8] ;
 wire \rbzero.traced_texa[9] ;
 wire \rbzero.vga_sync.vsync ;
 wire \rbzero.wall_hot[0] ;
 wire \rbzero.wall_hot[1] ;
 wire \rbzero.wall_tracer.mapX[10] ;
 wire \rbzero.wall_tracer.mapX[5] ;
 wire \rbzero.wall_tracer.mapX[6] ;
 wire \rbzero.wall_tracer.mapX[7] ;
 wire \rbzero.wall_tracer.mapX[8] ;
 wire \rbzero.wall_tracer.mapX[9] ;
 wire \rbzero.wall_tracer.mapY[10] ;
 wire \rbzero.wall_tracer.mapY[5] ;
 wire \rbzero.wall_tracer.mapY[6] ;
 wire \rbzero.wall_tracer.mapY[7] ;
 wire \rbzero.wall_tracer.mapY[8] ;
 wire \rbzero.wall_tracer.mapY[9] ;
 wire \rbzero.wall_tracer.rayAddendX[-1] ;
 wire \rbzero.wall_tracer.rayAddendX[-2] ;
 wire \rbzero.wall_tracer.rayAddendX[-3] ;
 wire \rbzero.wall_tracer.rayAddendX[-4] ;
 wire \rbzero.wall_tracer.rayAddendX[-5] ;
 wire \rbzero.wall_tracer.rayAddendX[-6] ;
 wire \rbzero.wall_tracer.rayAddendX[-7] ;
 wire \rbzero.wall_tracer.rayAddendX[-8] ;
 wire \rbzero.wall_tracer.rayAddendX[-9] ;
 wire \rbzero.wall_tracer.rayAddendX[0] ;
 wire \rbzero.wall_tracer.rayAddendX[10] ;
 wire \rbzero.wall_tracer.rayAddendX[1] ;
 wire \rbzero.wall_tracer.rayAddendX[2] ;
 wire \rbzero.wall_tracer.rayAddendX[3] ;
 wire \rbzero.wall_tracer.rayAddendX[4] ;
 wire \rbzero.wall_tracer.rayAddendX[5] ;
 wire \rbzero.wall_tracer.rayAddendX[6] ;
 wire \rbzero.wall_tracer.rayAddendX[7] ;
 wire \rbzero.wall_tracer.rayAddendX[8] ;
 wire \rbzero.wall_tracer.rayAddendX[9] ;
 wire \rbzero.wall_tracer.rayAddendY[-1] ;
 wire \rbzero.wall_tracer.rayAddendY[-2] ;
 wire \rbzero.wall_tracer.rayAddendY[-3] ;
 wire \rbzero.wall_tracer.rayAddendY[-4] ;
 wire \rbzero.wall_tracer.rayAddendY[-5] ;
 wire \rbzero.wall_tracer.rayAddendY[-6] ;
 wire \rbzero.wall_tracer.rayAddendY[-7] ;
 wire \rbzero.wall_tracer.rayAddendY[-8] ;
 wire \rbzero.wall_tracer.rayAddendY[-9] ;
 wire \rbzero.wall_tracer.rayAddendY[0] ;
 wire \rbzero.wall_tracer.rayAddendY[10] ;
 wire \rbzero.wall_tracer.rayAddendY[1] ;
 wire \rbzero.wall_tracer.rayAddendY[2] ;
 wire \rbzero.wall_tracer.rayAddendY[3] ;
 wire \rbzero.wall_tracer.rayAddendY[4] ;
 wire \rbzero.wall_tracer.rayAddendY[5] ;
 wire \rbzero.wall_tracer.rayAddendY[6] ;
 wire \rbzero.wall_tracer.rayAddendY[7] ;
 wire \rbzero.wall_tracer.rayAddendY[8] ;
 wire \rbzero.wall_tracer.rayAddendY[9] ;
 wire \rbzero.wall_tracer.rcp_sel[0] ;
 wire \rbzero.wall_tracer.rcp_sel[2] ;
 wire \rbzero.wall_tracer.stepDistX[-10] ;
 wire \rbzero.wall_tracer.stepDistX[-11] ;
 wire \rbzero.wall_tracer.stepDistX[-1] ;
 wire \rbzero.wall_tracer.stepDistX[-2] ;
 wire \rbzero.wall_tracer.stepDistX[-3] ;
 wire \rbzero.wall_tracer.stepDistX[-4] ;
 wire \rbzero.wall_tracer.stepDistX[-5] ;
 wire \rbzero.wall_tracer.stepDistX[-6] ;
 wire \rbzero.wall_tracer.stepDistX[-7] ;
 wire \rbzero.wall_tracer.stepDistX[-8] ;
 wire \rbzero.wall_tracer.stepDistX[-9] ;
 wire \rbzero.wall_tracer.stepDistX[0] ;
 wire \rbzero.wall_tracer.stepDistX[10] ;
 wire \rbzero.wall_tracer.stepDistX[1] ;
 wire \rbzero.wall_tracer.stepDistX[2] ;
 wire \rbzero.wall_tracer.stepDistX[3] ;
 wire \rbzero.wall_tracer.stepDistX[4] ;
 wire \rbzero.wall_tracer.stepDistX[5] ;
 wire \rbzero.wall_tracer.stepDistX[6] ;
 wire \rbzero.wall_tracer.stepDistX[7] ;
 wire \rbzero.wall_tracer.stepDistX[8] ;
 wire \rbzero.wall_tracer.stepDistX[9] ;
 wire \rbzero.wall_tracer.stepDistY[-10] ;
 wire \rbzero.wall_tracer.stepDistY[-11] ;
 wire \rbzero.wall_tracer.stepDistY[-1] ;
 wire \rbzero.wall_tracer.stepDistY[-2] ;
 wire \rbzero.wall_tracer.stepDistY[-3] ;
 wire \rbzero.wall_tracer.stepDistY[-4] ;
 wire \rbzero.wall_tracer.stepDistY[-5] ;
 wire \rbzero.wall_tracer.stepDistY[-6] ;
 wire \rbzero.wall_tracer.stepDistY[-7] ;
 wire \rbzero.wall_tracer.stepDistY[-8] ;
 wire \rbzero.wall_tracer.stepDistY[-9] ;
 wire \rbzero.wall_tracer.stepDistY[0] ;
 wire \rbzero.wall_tracer.stepDistY[10] ;
 wire \rbzero.wall_tracer.stepDistY[1] ;
 wire \rbzero.wall_tracer.stepDistY[2] ;
 wire \rbzero.wall_tracer.stepDistY[3] ;
 wire \rbzero.wall_tracer.stepDistY[4] ;
 wire \rbzero.wall_tracer.stepDistY[5] ;
 wire \rbzero.wall_tracer.stepDistY[6] ;
 wire \rbzero.wall_tracer.stepDistY[7] ;
 wire \rbzero.wall_tracer.stepDistY[8] ;
 wire \rbzero.wall_tracer.stepDistY[9] ;
 wire \rbzero.wall_tracer.trackDistX[-10] ;
 wire \rbzero.wall_tracer.trackDistX[-11] ;
 wire \rbzero.wall_tracer.trackDistX[-1] ;
 wire \rbzero.wall_tracer.trackDistX[-2] ;
 wire \rbzero.wall_tracer.trackDistX[-3] ;
 wire \rbzero.wall_tracer.trackDistX[-4] ;
 wire \rbzero.wall_tracer.trackDistX[-5] ;
 wire \rbzero.wall_tracer.trackDistX[-6] ;
 wire \rbzero.wall_tracer.trackDistX[-7] ;
 wire \rbzero.wall_tracer.trackDistX[-8] ;
 wire \rbzero.wall_tracer.trackDistX[-9] ;
 wire \rbzero.wall_tracer.trackDistX[0] ;
 wire \rbzero.wall_tracer.trackDistX[10] ;
 wire \rbzero.wall_tracer.trackDistX[1] ;
 wire \rbzero.wall_tracer.trackDistX[2] ;
 wire \rbzero.wall_tracer.trackDistX[3] ;
 wire \rbzero.wall_tracer.trackDistX[4] ;
 wire \rbzero.wall_tracer.trackDistX[5] ;
 wire \rbzero.wall_tracer.trackDistX[6] ;
 wire \rbzero.wall_tracer.trackDistX[7] ;
 wire \rbzero.wall_tracer.trackDistX[8] ;
 wire \rbzero.wall_tracer.trackDistX[9] ;
 wire \rbzero.wall_tracer.trackDistY[-10] ;
 wire \rbzero.wall_tracer.trackDistY[-11] ;
 wire \rbzero.wall_tracer.trackDistY[-1] ;
 wire \rbzero.wall_tracer.trackDistY[-2] ;
 wire \rbzero.wall_tracer.trackDistY[-3] ;
 wire \rbzero.wall_tracer.trackDistY[-4] ;
 wire \rbzero.wall_tracer.trackDistY[-5] ;
 wire \rbzero.wall_tracer.trackDistY[-6] ;
 wire \rbzero.wall_tracer.trackDistY[-7] ;
 wire \rbzero.wall_tracer.trackDistY[-8] ;
 wire \rbzero.wall_tracer.trackDistY[-9] ;
 wire \rbzero.wall_tracer.trackDistY[0] ;
 wire \rbzero.wall_tracer.trackDistY[10] ;
 wire \rbzero.wall_tracer.trackDistY[1] ;
 wire \rbzero.wall_tracer.trackDistY[2] ;
 wire \rbzero.wall_tracer.trackDistY[3] ;
 wire \rbzero.wall_tracer.trackDistY[4] ;
 wire \rbzero.wall_tracer.trackDistY[5] ;
 wire \rbzero.wall_tracer.trackDistY[6] ;
 wire \rbzero.wall_tracer.trackDistY[7] ;
 wire \rbzero.wall_tracer.trackDistY[8] ;
 wire \rbzero.wall_tracer.trackDistY[9] ;
 wire \rbzero.wall_tracer.visualWallDist[-10] ;
 wire \rbzero.wall_tracer.visualWallDist[-11] ;
 wire \rbzero.wall_tracer.visualWallDist[-1] ;
 wire \rbzero.wall_tracer.visualWallDist[-2] ;
 wire \rbzero.wall_tracer.visualWallDist[-3] ;
 wire \rbzero.wall_tracer.visualWallDist[-4] ;
 wire \rbzero.wall_tracer.visualWallDist[-5] ;
 wire \rbzero.wall_tracer.visualWallDist[-6] ;
 wire \rbzero.wall_tracer.visualWallDist[-7] ;
 wire \rbzero.wall_tracer.visualWallDist[-8] ;
 wire \rbzero.wall_tracer.visualWallDist[-9] ;
 wire \rbzero.wall_tracer.visualWallDist[0] ;
 wire \rbzero.wall_tracer.visualWallDist[10] ;
 wire \rbzero.wall_tracer.visualWallDist[1] ;
 wire \rbzero.wall_tracer.visualWallDist[2] ;
 wire \rbzero.wall_tracer.visualWallDist[3] ;
 wire \rbzero.wall_tracer.visualWallDist[4] ;
 wire \rbzero.wall_tracer.visualWallDist[5] ;
 wire \rbzero.wall_tracer.visualWallDist[6] ;
 wire \rbzero.wall_tracer.visualWallDist[7] ;
 wire \rbzero.wall_tracer.visualWallDist[8] ;
 wire \rbzero.wall_tracer.visualWallDist[9] ;
 wire \reg_gpout[0] ;
 wire \reg_gpout[1] ;
 wire \reg_gpout[2] ;
 wire \reg_gpout[3] ;
 wire \reg_gpout[4] ;
 wire \reg_gpout[5] ;
 wire reg_hsync;
 wire \reg_rgb[14] ;
 wire \reg_rgb[15] ;
 wire \reg_rgb[22] ;
 wire \reg_rgb[23] ;
 wire \reg_rgb[6] ;
 wire \reg_rgb[7] ;
 wire reg_vsync;
 wire net94;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net127;
 wire net74;
 wire net75;
 wire net126;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_9_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_52_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_62_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_65_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_67_i_clk;
 wire clknet_leaf_68_i_clk;
 wire clknet_leaf_69_i_clk;
 wire clknet_leaf_70_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_72_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_79_i_clk;
 wire clknet_leaf_80_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_82_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_86_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_90_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_94_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_leaf_96_i_clk;
 wire clknet_leaf_97_i_clk;
 wire clknet_leaf_98_i_clk;
 wire clknet_leaf_99_i_clk;
 wire clknet_leaf_100_i_clk;
 wire clknet_0_i_clk;
 wire clknet_1_0_0_i_clk;
 wire clknet_1_0_1_i_clk;
 wire clknet_1_1_0_i_clk;
 wire clknet_1_1_1_i_clk;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_3_0_i_clk;
 wire clknet_3_0_0_i_clk;
 wire clknet_3_1_0_i_clk;
 wire clknet_3_2_0_i_clk;
 wire clknet_3_3_0_i_clk;
 wire clknet_3_4_0_i_clk;
 wire clknet_3_5_0_i_clk;
 wire clknet_3_6_0_i_clk;
 wire clknet_3_7_0_i_clk;
 wire clknet_opt_1_0_i_clk;
 wire clknet_opt_2_0_i_clk;
 wire clknet_opt_3_0_i_clk;
 wire clknet_opt_4_0_i_clk;
 wire clknet_0__05820_;
 wire clknet_1_0__leaf__05820_;
 wire clknet_1_1__leaf__05820_;
 wire clknet_0__05700_;
 wire clknet_1_0__leaf__05700_;
 wire clknet_1_1__leaf__05700_;
 wire clknet_0__04634_;
 wire clknet_1_0__leaf__04634_;
 wire clknet_1_1__leaf__04634_;
 wire clknet_0__05993_;
 wire clknet_1_0__leaf__05993_;
 wire clknet_1_1__leaf__05993_;
 wire clknet_0__03808_;
 wire clknet_1_0__leaf__03808_;
 wire clknet_1_1__leaf__03808_;
 wire clknet_0__03807_;
 wire clknet_1_0__leaf__03807_;
 wire clknet_1_1__leaf__03807_;
 wire clknet_0__03796_;
 wire clknet_1_0__leaf__03796_;
 wire clknet_1_1__leaf__03796_;
 wire clknet_0__03806_;
 wire clknet_1_0__leaf__03806_;
 wire clknet_1_1__leaf__03806_;
 wire clknet_0__03805_;
 wire clknet_1_0__leaf__03805_;
 wire clknet_1_1__leaf__03805_;
 wire clknet_0__03804_;
 wire clknet_1_0__leaf__03804_;
 wire clknet_1_1__leaf__03804_;
 wire clknet_0__03803_;
 wire clknet_1_0__leaf__03803_;
 wire clknet_1_1__leaf__03803_;
 wire clknet_0__03802_;
 wire clknet_1_0__leaf__03802_;
 wire clknet_1_1__leaf__03802_;
 wire clknet_0__03801_;
 wire clknet_1_0__leaf__03801_;
 wire clknet_1_1__leaf__03801_;
 wire clknet_0__03800_;
 wire clknet_1_0__leaf__03800_;
 wire clknet_1_1__leaf__03800_;
 wire clknet_0__03799_;
 wire clknet_1_0__leaf__03799_;
 wire clknet_1_1__leaf__03799_;
 wire clknet_0__03798_;
 wire clknet_1_0__leaf__03798_;
 wire clknet_1_1__leaf__03798_;
 wire clknet_0__03797_;
 wire clknet_1_0__leaf__03797_;
 wire clknet_1_1__leaf__03797_;
 wire clknet_0__03785_;
 wire clknet_1_0__leaf__03785_;
 wire clknet_1_1__leaf__03785_;
 wire clknet_0__03795_;
 wire clknet_1_0__leaf__03795_;
 wire clknet_1_1__leaf__03795_;
 wire clknet_0__03794_;
 wire clknet_1_0__leaf__03794_;
 wire clknet_1_1__leaf__03794_;
 wire clknet_0__03793_;
 wire clknet_1_0__leaf__03793_;
 wire clknet_1_1__leaf__03793_;
 wire clknet_0__03792_;
 wire clknet_1_0__leaf__03792_;
 wire clknet_1_1__leaf__03792_;
 wire clknet_0__03791_;
 wire clknet_1_0__leaf__03791_;
 wire clknet_1_1__leaf__03791_;
 wire clknet_0__03790_;
 wire clknet_1_0__leaf__03790_;
 wire clknet_1_1__leaf__03790_;
 wire clknet_0__03789_;
 wire clknet_1_0__leaf__03789_;
 wire clknet_1_1__leaf__03789_;
 wire clknet_0__03788_;
 wire clknet_1_0__leaf__03788_;
 wire clknet_1_1__leaf__03788_;
 wire clknet_0__03787_;
 wire clknet_1_0__leaf__03787_;
 wire clknet_1_1__leaf__03787_;
 wire clknet_0__03786_;
 wire clknet_1_0__leaf__03786_;
 wire clknet_1_1__leaf__03786_;
 wire clknet_0__03464_;
 wire clknet_1_0__leaf__03464_;
 wire clknet_1_1__leaf__03464_;
 wire clknet_0__03784_;
 wire clknet_1_0__leaf__03784_;
 wire clknet_1_1__leaf__03784_;
 wire clknet_0__03783_;
 wire clknet_1_0__leaf__03783_;
 wire clknet_1_1__leaf__03783_;
 wire clknet_0__03782_;
 wire clknet_1_0__leaf__03782_;
 wire clknet_1_1__leaf__03782_;
 wire clknet_0__03781_;
 wire clknet_1_0__leaf__03781_;
 wire clknet_1_1__leaf__03781_;
 wire clknet_0__03780_;
 wire clknet_1_0__leaf__03780_;
 wire clknet_1_1__leaf__03780_;
 wire clknet_0__03779_;
 wire clknet_1_0__leaf__03779_;
 wire clknet_1_1__leaf__03779_;
 wire clknet_0__03778_;
 wire clknet_1_0__leaf__03778_;
 wire clknet_1_1__leaf__03778_;
 wire clknet_0__03777_;
 wire clknet_1_0__leaf__03777_;
 wire clknet_1_1__leaf__03777_;
 wire clknet_0__03776_;
 wire clknet_1_0__leaf__03776_;
 wire clknet_1_1__leaf__03776_;
 wire clknet_0__03465_;
 wire clknet_1_0__leaf__03465_;
 wire clknet_1_1__leaf__03465_;
 wire clknet_0__03457_;
 wire clknet_1_0__leaf__03457_;
 wire clknet_1_1__leaf__03457_;
 wire clknet_0__03463_;
 wire clknet_1_0__leaf__03463_;
 wire clknet_1_1__leaf__03463_;
 wire clknet_0__03462_;
 wire clknet_1_0__leaf__03462_;
 wire clknet_1_1__leaf__03462_;
 wire clknet_0__03461_;
 wire clknet_1_0__leaf__03461_;
 wire clknet_1_1__leaf__03461_;
 wire clknet_0__03460_;
 wire clknet_1_0__leaf__03460_;
 wire clknet_1_1__leaf__03460_;
 wire clknet_0__03459_;
 wire clknet_1_0__leaf__03459_;
 wire clknet_1_1__leaf__03459_;
 wire clknet_0__03458_;
 wire clknet_1_0__leaf__03458_;
 wire clknet_1_1__leaf__03458_;
 wire clknet_0__05938_;
 wire clknet_1_0__leaf__05938_;
 wire clknet_1_1__leaf__05938_;
 wire clknet_0__05879_;
 wire clknet_1_0__leaf__05879_;
 wire clknet_1_1__leaf__05879_;
 wire clknet_0__05761_;
 wire clknet_1_0__leaf__05761_;
 wire clknet_1_1__leaf__05761_;
 wire net73;
 wire net511;
 wire net512;

 sky130_fd_sc_hd__buf_4 _10388_ (.A(\gpout0.hpos[0] ),
    .X(_03969_));
 sky130_fd_sc_hd__clkbuf_4 _10389_ (.A(_03969_),
    .X(_03970_));
 sky130_fd_sc_hd__buf_4 _10390_ (.A(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__buf_4 _10391_ (.A(\gpout0.hpos[7] ),
    .X(_03972_));
 sky130_fd_sc_hd__clkbuf_4 _10392_ (.A(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__xor2_4 _10393_ (.A(net47),
    .B(net48),
    .X(_03974_));
 sky130_fd_sc_hd__clkbuf_4 _10394_ (.A(\gpout0.hpos[8] ),
    .X(_03975_));
 sky130_fd_sc_hd__inv_2 _10395_ (.A(\gpout0.hpos[9] ),
    .Y(_03976_));
 sky130_fd_sc_hd__nor2_1 _10396_ (.A(_03975_),
    .B(_03976_),
    .Y(_03977_));
 sky130_fd_sc_hd__and4_2 _10397_ (.A(_03971_),
    .B(_03973_),
    .C(_03974_),
    .D(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__buf_4 _10398_ (.A(_03978_),
    .X(_03979_));
 sky130_fd_sc_hd__clkbuf_4 _10399_ (.A(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__mux2_1 _10400_ (.A0(\rbzero.tex_r1[63] ),
    .A1(net49),
    .S(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__clkbuf_1 _10401_ (.A(_03981_),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _10402_ (.A0(\rbzero.tex_r1[62] ),
    .A1(\rbzero.tex_r1[63] ),
    .S(_03980_),
    .X(_03982_));
 sky130_fd_sc_hd__clkbuf_1 _10403_ (.A(_03982_),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _10404_ (.A0(\rbzero.tex_r1[61] ),
    .A1(\rbzero.tex_r1[62] ),
    .S(_03980_),
    .X(_03983_));
 sky130_fd_sc_hd__clkbuf_1 _10405_ (.A(_03983_),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _10406_ (.A0(\rbzero.tex_r1[60] ),
    .A1(\rbzero.tex_r1[61] ),
    .S(_03980_),
    .X(_03984_));
 sky130_fd_sc_hd__clkbuf_1 _10407_ (.A(_03984_),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _10408_ (.A0(\rbzero.tex_r1[59] ),
    .A1(\rbzero.tex_r1[60] ),
    .S(_03980_),
    .X(_03985_));
 sky130_fd_sc_hd__clkbuf_1 _10409_ (.A(_03985_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _10410_ (.A0(\rbzero.tex_r1[58] ),
    .A1(\rbzero.tex_r1[59] ),
    .S(_03980_),
    .X(_03986_));
 sky130_fd_sc_hd__clkbuf_1 _10411_ (.A(_03986_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _10412_ (.A0(\rbzero.tex_r1[57] ),
    .A1(\rbzero.tex_r1[58] ),
    .S(_03980_),
    .X(_03987_));
 sky130_fd_sc_hd__clkbuf_1 _10413_ (.A(_03987_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _10414_ (.A0(\rbzero.tex_r1[56] ),
    .A1(\rbzero.tex_r1[57] ),
    .S(_03980_),
    .X(_03988_));
 sky130_fd_sc_hd__clkbuf_1 _10415_ (.A(_03988_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _10416_ (.A0(\rbzero.tex_r1[55] ),
    .A1(\rbzero.tex_r1[56] ),
    .S(_03980_),
    .X(_03989_));
 sky130_fd_sc_hd__clkbuf_1 _10417_ (.A(_03989_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _10418_ (.A0(\rbzero.tex_r1[54] ),
    .A1(\rbzero.tex_r1[55] ),
    .S(_03980_),
    .X(_03990_));
 sky130_fd_sc_hd__clkbuf_1 _10419_ (.A(_03990_),
    .X(_01588_));
 sky130_fd_sc_hd__clkbuf_4 _10420_ (.A(_03979_),
    .X(_03991_));
 sky130_fd_sc_hd__mux2_1 _10421_ (.A0(\rbzero.tex_r1[53] ),
    .A1(\rbzero.tex_r1[54] ),
    .S(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__clkbuf_1 _10422_ (.A(_03992_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _10423_ (.A0(\rbzero.tex_r1[52] ),
    .A1(\rbzero.tex_r1[53] ),
    .S(_03991_),
    .X(_03993_));
 sky130_fd_sc_hd__clkbuf_1 _10424_ (.A(_03993_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _10425_ (.A0(\rbzero.tex_r1[51] ),
    .A1(\rbzero.tex_r1[52] ),
    .S(_03991_),
    .X(_03994_));
 sky130_fd_sc_hd__clkbuf_1 _10426_ (.A(_03994_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _10427_ (.A0(\rbzero.tex_r1[50] ),
    .A1(\rbzero.tex_r1[51] ),
    .S(_03991_),
    .X(_03995_));
 sky130_fd_sc_hd__clkbuf_1 _10428_ (.A(_03995_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _10429_ (.A0(\rbzero.tex_r1[49] ),
    .A1(\rbzero.tex_r1[50] ),
    .S(_03991_),
    .X(_03996_));
 sky130_fd_sc_hd__clkbuf_1 _10430_ (.A(_03996_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _10431_ (.A0(\rbzero.tex_r1[48] ),
    .A1(\rbzero.tex_r1[49] ),
    .S(_03991_),
    .X(_03997_));
 sky130_fd_sc_hd__clkbuf_1 _10432_ (.A(_03997_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _10433_ (.A0(\rbzero.tex_r1[47] ),
    .A1(\rbzero.tex_r1[48] ),
    .S(_03991_),
    .X(_03998_));
 sky130_fd_sc_hd__clkbuf_1 _10434_ (.A(_03998_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _10435_ (.A0(\rbzero.tex_r1[46] ),
    .A1(\rbzero.tex_r1[47] ),
    .S(_03991_),
    .X(_03999_));
 sky130_fd_sc_hd__clkbuf_1 _10436_ (.A(_03999_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _10437_ (.A0(\rbzero.tex_r1[45] ),
    .A1(\rbzero.tex_r1[46] ),
    .S(_03991_),
    .X(_04000_));
 sky130_fd_sc_hd__clkbuf_1 _10438_ (.A(_04000_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _10439_ (.A0(\rbzero.tex_r1[44] ),
    .A1(\rbzero.tex_r1[45] ),
    .S(_03991_),
    .X(_04001_));
 sky130_fd_sc_hd__clkbuf_1 _10440_ (.A(_04001_),
    .X(_01578_));
 sky130_fd_sc_hd__clkbuf_4 _10441_ (.A(_03979_),
    .X(_04002_));
 sky130_fd_sc_hd__mux2_1 _10442_ (.A0(\rbzero.tex_r1[43] ),
    .A1(\rbzero.tex_r1[44] ),
    .S(_04002_),
    .X(_04003_));
 sky130_fd_sc_hd__clkbuf_1 _10443_ (.A(_04003_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _10444_ (.A0(\rbzero.tex_r1[42] ),
    .A1(\rbzero.tex_r1[43] ),
    .S(_04002_),
    .X(_04004_));
 sky130_fd_sc_hd__clkbuf_1 _10445_ (.A(_04004_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _10446_ (.A0(\rbzero.tex_r1[41] ),
    .A1(\rbzero.tex_r1[42] ),
    .S(_04002_),
    .X(_04005_));
 sky130_fd_sc_hd__clkbuf_1 _10447_ (.A(_04005_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _10448_ (.A0(\rbzero.tex_r1[40] ),
    .A1(\rbzero.tex_r1[41] ),
    .S(_04002_),
    .X(_04006_));
 sky130_fd_sc_hd__clkbuf_1 _10449_ (.A(_04006_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _10450_ (.A0(\rbzero.tex_r1[39] ),
    .A1(net73),
    .S(_04002_),
    .X(_04007_));
 sky130_fd_sc_hd__clkbuf_1 _10451_ (.A(_04007_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _10452_ (.A0(\rbzero.tex_r1[38] ),
    .A1(\rbzero.tex_r1[39] ),
    .S(_04002_),
    .X(_04008_));
 sky130_fd_sc_hd__clkbuf_1 _10453_ (.A(_04008_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _10454_ (.A0(\rbzero.tex_r1[37] ),
    .A1(\rbzero.tex_r1[38] ),
    .S(_04002_),
    .X(_04009_));
 sky130_fd_sc_hd__clkbuf_1 _10455_ (.A(_04009_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _10456_ (.A0(\rbzero.tex_r1[36] ),
    .A1(\rbzero.tex_r1[37] ),
    .S(_04002_),
    .X(_04010_));
 sky130_fd_sc_hd__clkbuf_1 _10457_ (.A(_04010_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _10458_ (.A0(\rbzero.tex_r1[35] ),
    .A1(\rbzero.tex_r1[36] ),
    .S(_04002_),
    .X(_04011_));
 sky130_fd_sc_hd__clkbuf_1 _10459_ (.A(_04011_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(\rbzero.tex_r1[34] ),
    .A1(\rbzero.tex_r1[35] ),
    .S(_04002_),
    .X(_04012_));
 sky130_fd_sc_hd__clkbuf_1 _10461_ (.A(_04012_),
    .X(_01568_));
 sky130_fd_sc_hd__clkbuf_4 _10462_ (.A(_03979_),
    .X(_04013_));
 sky130_fd_sc_hd__mux2_1 _10463_ (.A0(\rbzero.tex_r1[33] ),
    .A1(\rbzero.tex_r1[34] ),
    .S(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__clkbuf_1 _10464_ (.A(_04014_),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _10465_ (.A0(\rbzero.tex_r1[32] ),
    .A1(\rbzero.tex_r1[33] ),
    .S(_04013_),
    .X(_04015_));
 sky130_fd_sc_hd__clkbuf_1 _10466_ (.A(_04015_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _10467_ (.A0(\rbzero.tex_r1[31] ),
    .A1(\rbzero.tex_r1[32] ),
    .S(_04013_),
    .X(_04016_));
 sky130_fd_sc_hd__clkbuf_1 _10468_ (.A(_04016_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _10469_ (.A0(\rbzero.tex_r1[30] ),
    .A1(\rbzero.tex_r1[31] ),
    .S(_04013_),
    .X(_04017_));
 sky130_fd_sc_hd__clkbuf_1 _10470_ (.A(_04017_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _10471_ (.A0(\rbzero.tex_r1[29] ),
    .A1(\rbzero.tex_r1[30] ),
    .S(_04013_),
    .X(_04018_));
 sky130_fd_sc_hd__clkbuf_1 _10472_ (.A(_04018_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _10473_ (.A0(\rbzero.tex_r1[28] ),
    .A1(\rbzero.tex_r1[29] ),
    .S(_04013_),
    .X(_04019_));
 sky130_fd_sc_hd__clkbuf_1 _10474_ (.A(_04019_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _10475_ (.A0(\rbzero.tex_r1[27] ),
    .A1(\rbzero.tex_r1[28] ),
    .S(_04013_),
    .X(_04020_));
 sky130_fd_sc_hd__clkbuf_1 _10476_ (.A(_04020_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(\rbzero.tex_r1[26] ),
    .A1(\rbzero.tex_r1[27] ),
    .S(_04013_),
    .X(_04021_));
 sky130_fd_sc_hd__clkbuf_1 _10478_ (.A(_04021_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(\rbzero.tex_r1[25] ),
    .A1(\rbzero.tex_r1[26] ),
    .S(_04013_),
    .X(_04022_));
 sky130_fd_sc_hd__clkbuf_1 _10480_ (.A(_04022_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _10481_ (.A0(\rbzero.tex_r1[24] ),
    .A1(\rbzero.tex_r1[25] ),
    .S(_04013_),
    .X(_04023_));
 sky130_fd_sc_hd__clkbuf_1 _10482_ (.A(_04023_),
    .X(_01558_));
 sky130_fd_sc_hd__clkbuf_4 _10483_ (.A(_03979_),
    .X(_04024_));
 sky130_fd_sc_hd__mux2_1 _10484_ (.A0(\rbzero.tex_r1[23] ),
    .A1(\rbzero.tex_r1[24] ),
    .S(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__clkbuf_1 _10485_ (.A(_04025_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _10486_ (.A0(\rbzero.tex_r1[22] ),
    .A1(\rbzero.tex_r1[23] ),
    .S(_04024_),
    .X(_04026_));
 sky130_fd_sc_hd__clkbuf_1 _10487_ (.A(_04026_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _10488_ (.A0(\rbzero.tex_r1[21] ),
    .A1(\rbzero.tex_r1[22] ),
    .S(_04024_),
    .X(_04027_));
 sky130_fd_sc_hd__clkbuf_1 _10489_ (.A(_04027_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _10490_ (.A0(\rbzero.tex_r1[20] ),
    .A1(\rbzero.tex_r1[21] ),
    .S(_04024_),
    .X(_04028_));
 sky130_fd_sc_hd__clkbuf_1 _10491_ (.A(_04028_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _10492_ (.A0(\rbzero.tex_r1[19] ),
    .A1(\rbzero.tex_r1[20] ),
    .S(_04024_),
    .X(_04029_));
 sky130_fd_sc_hd__clkbuf_1 _10493_ (.A(_04029_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _10494_ (.A0(\rbzero.tex_r1[18] ),
    .A1(\rbzero.tex_r1[19] ),
    .S(_04024_),
    .X(_04030_));
 sky130_fd_sc_hd__clkbuf_1 _10495_ (.A(_04030_),
    .X(_01552_));
 sky130_fd_sc_hd__mux2_1 _10496_ (.A0(\rbzero.tex_r1[17] ),
    .A1(\rbzero.tex_r1[18] ),
    .S(_04024_),
    .X(_04031_));
 sky130_fd_sc_hd__clkbuf_1 _10497_ (.A(_04031_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _10498_ (.A0(\rbzero.tex_r1[16] ),
    .A1(\rbzero.tex_r1[17] ),
    .S(_04024_),
    .X(_04032_));
 sky130_fd_sc_hd__clkbuf_1 _10499_ (.A(_04032_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _10500_ (.A0(\rbzero.tex_r1[15] ),
    .A1(\rbzero.tex_r1[16] ),
    .S(_04024_),
    .X(_04033_));
 sky130_fd_sc_hd__clkbuf_1 _10501_ (.A(_04033_),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _10502_ (.A0(\rbzero.tex_r1[14] ),
    .A1(\rbzero.tex_r1[15] ),
    .S(_04024_),
    .X(_04034_));
 sky130_fd_sc_hd__clkbuf_1 _10503_ (.A(_04034_),
    .X(_01548_));
 sky130_fd_sc_hd__clkbuf_4 _10504_ (.A(_03979_),
    .X(_04035_));
 sky130_fd_sc_hd__mux2_1 _10505_ (.A0(\rbzero.tex_r1[13] ),
    .A1(\rbzero.tex_r1[14] ),
    .S(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__clkbuf_1 _10506_ (.A(_04036_),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _10507_ (.A0(\rbzero.tex_r1[12] ),
    .A1(\rbzero.tex_r1[13] ),
    .S(_04035_),
    .X(_04037_));
 sky130_fd_sc_hd__clkbuf_1 _10508_ (.A(_04037_),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _10509_ (.A0(\rbzero.tex_r1[11] ),
    .A1(\rbzero.tex_r1[12] ),
    .S(_04035_),
    .X(_04038_));
 sky130_fd_sc_hd__clkbuf_1 _10510_ (.A(_04038_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(\rbzero.tex_r1[10] ),
    .A1(\rbzero.tex_r1[11] ),
    .S(_04035_),
    .X(_04039_));
 sky130_fd_sc_hd__clkbuf_1 _10512_ (.A(_04039_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _10513_ (.A0(\rbzero.tex_r1[9] ),
    .A1(\rbzero.tex_r1[10] ),
    .S(_04035_),
    .X(_04040_));
 sky130_fd_sc_hd__clkbuf_1 _10514_ (.A(_04040_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(\rbzero.tex_r1[8] ),
    .A1(\rbzero.tex_r1[9] ),
    .S(_04035_),
    .X(_04041_));
 sky130_fd_sc_hd__clkbuf_1 _10516_ (.A(_04041_),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(\rbzero.tex_r1[7] ),
    .A1(\rbzero.tex_r1[8] ),
    .S(_04035_),
    .X(_04042_));
 sky130_fd_sc_hd__clkbuf_1 _10518_ (.A(_04042_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _10519_ (.A0(\rbzero.tex_r1[6] ),
    .A1(\rbzero.tex_r1[7] ),
    .S(_04035_),
    .X(_04043_));
 sky130_fd_sc_hd__clkbuf_1 _10520_ (.A(_04043_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(\rbzero.tex_r1[5] ),
    .A1(\rbzero.tex_r1[6] ),
    .S(_04035_),
    .X(_04044_));
 sky130_fd_sc_hd__clkbuf_1 _10522_ (.A(_04044_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _10523_ (.A0(\rbzero.tex_r1[4] ),
    .A1(\rbzero.tex_r1[5] ),
    .S(_04035_),
    .X(_04045_));
 sky130_fd_sc_hd__clkbuf_1 _10524_ (.A(_04045_),
    .X(_01538_));
 sky130_fd_sc_hd__clkbuf_4 _10525_ (.A(_03979_),
    .X(_04046_));
 sky130_fd_sc_hd__mux2_1 _10526_ (.A0(\rbzero.tex_r1[3] ),
    .A1(\rbzero.tex_r1[4] ),
    .S(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__clkbuf_1 _10527_ (.A(_04047_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _10528_ (.A0(\rbzero.tex_r1[2] ),
    .A1(\rbzero.tex_r1[3] ),
    .S(_04046_),
    .X(_04048_));
 sky130_fd_sc_hd__clkbuf_1 _10529_ (.A(_04048_),
    .X(_01536_));
 sky130_fd_sc_hd__mux2_1 _10530_ (.A0(\rbzero.tex_r1[1] ),
    .A1(\rbzero.tex_r1[2] ),
    .S(_04046_),
    .X(_04049_));
 sky130_fd_sc_hd__clkbuf_1 _10531_ (.A(_04049_),
    .X(_01535_));
 sky130_fd_sc_hd__mux2_1 _10532_ (.A0(\rbzero.tex_r1[0] ),
    .A1(\rbzero.tex_r1[1] ),
    .S(_04046_),
    .X(_04050_));
 sky130_fd_sc_hd__clkbuf_1 _10533_ (.A(_04050_),
    .X(_01534_));
 sky130_fd_sc_hd__inv_2 _10534_ (.A(_03973_),
    .Y(_04051_));
 sky130_fd_sc_hd__clkinv_4 _10535_ (.A(_03974_),
    .Y(_04052_));
 sky130_fd_sc_hd__or4b_4 _10536_ (.A(_03971_),
    .B(_04051_),
    .C(_04052_),
    .D_N(_03977_),
    .X(_04053_));
 sky130_fd_sc_hd__buf_4 _10537_ (.A(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__clkbuf_4 _10538_ (.A(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__mux2_1 _10539_ (.A0(net49),
    .A1(\rbzero.tex_r0[63] ),
    .S(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__clkbuf_1 _10540_ (.A(_04056_),
    .X(_01533_));
 sky130_fd_sc_hd__mux2_1 _10541_ (.A0(\rbzero.tex_r0[63] ),
    .A1(\rbzero.tex_r0[62] ),
    .S(_04055_),
    .X(_04057_));
 sky130_fd_sc_hd__clkbuf_1 _10542_ (.A(_04057_),
    .X(_01532_));
 sky130_fd_sc_hd__mux2_1 _10543_ (.A0(\rbzero.tex_r0[62] ),
    .A1(\rbzero.tex_r0[61] ),
    .S(_04055_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_1 _10544_ (.A(_04058_),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _10545_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_04055_),
    .X(_04059_));
 sky130_fd_sc_hd__clkbuf_1 _10546_ (.A(_04059_),
    .X(_01530_));
 sky130_fd_sc_hd__mux2_1 _10547_ (.A0(\rbzero.tex_r0[60] ),
    .A1(\rbzero.tex_r0[59] ),
    .S(_04055_),
    .X(_04060_));
 sky130_fd_sc_hd__clkbuf_1 _10548_ (.A(_04060_),
    .X(_01529_));
 sky130_fd_sc_hd__mux2_1 _10549_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_04055_),
    .X(_04061_));
 sky130_fd_sc_hd__clkbuf_1 _10550_ (.A(_04061_),
    .X(_01528_));
 sky130_fd_sc_hd__mux2_1 _10551_ (.A0(\rbzero.tex_r0[58] ),
    .A1(\rbzero.tex_r0[57] ),
    .S(_04055_),
    .X(_04062_));
 sky130_fd_sc_hd__clkbuf_1 _10552_ (.A(_04062_),
    .X(_01527_));
 sky130_fd_sc_hd__mux2_1 _10553_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_04055_),
    .X(_04063_));
 sky130_fd_sc_hd__clkbuf_1 _10554_ (.A(_04063_),
    .X(_01526_));
 sky130_fd_sc_hd__mux2_1 _10555_ (.A0(\rbzero.tex_r0[56] ),
    .A1(\rbzero.tex_r0[55] ),
    .S(_04055_),
    .X(_04064_));
 sky130_fd_sc_hd__clkbuf_1 _10556_ (.A(_04064_),
    .X(_01525_));
 sky130_fd_sc_hd__mux2_1 _10557_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_04055_),
    .X(_04065_));
 sky130_fd_sc_hd__clkbuf_1 _10558_ (.A(_04065_),
    .X(_01524_));
 sky130_fd_sc_hd__clkbuf_4 _10559_ (.A(_04054_),
    .X(_04066_));
 sky130_fd_sc_hd__mux2_1 _10560_ (.A0(\rbzero.tex_r0[54] ),
    .A1(\rbzero.tex_r0[53] ),
    .S(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__clkbuf_1 _10561_ (.A(_04067_),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _10562_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_04066_),
    .X(_04068_));
 sky130_fd_sc_hd__clkbuf_1 _10563_ (.A(_04068_),
    .X(_01522_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(\rbzero.tex_r0[52] ),
    .A1(\rbzero.tex_r0[51] ),
    .S(_04066_),
    .X(_04069_));
 sky130_fd_sc_hd__clkbuf_1 _10565_ (.A(_04069_),
    .X(_01521_));
 sky130_fd_sc_hd__mux2_1 _10566_ (.A0(\rbzero.tex_r0[51] ),
    .A1(\rbzero.tex_r0[50] ),
    .S(_04066_),
    .X(_04070_));
 sky130_fd_sc_hd__clkbuf_1 _10567_ (.A(_04070_),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _10568_ (.A0(\rbzero.tex_r0[50] ),
    .A1(\rbzero.tex_r0[49] ),
    .S(_04066_),
    .X(_04071_));
 sky130_fd_sc_hd__clkbuf_1 _10569_ (.A(_04071_),
    .X(_01519_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_04066_),
    .X(_04072_));
 sky130_fd_sc_hd__clkbuf_1 _10571_ (.A(_04072_),
    .X(_01518_));
 sky130_fd_sc_hd__mux2_1 _10572_ (.A0(\rbzero.tex_r0[48] ),
    .A1(\rbzero.tex_r0[47] ),
    .S(_04066_),
    .X(_04073_));
 sky130_fd_sc_hd__clkbuf_1 _10573_ (.A(_04073_),
    .X(_01517_));
 sky130_fd_sc_hd__mux2_1 _10574_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_04066_),
    .X(_04074_));
 sky130_fd_sc_hd__clkbuf_1 _10575_ (.A(_04074_),
    .X(_01516_));
 sky130_fd_sc_hd__mux2_1 _10576_ (.A0(\rbzero.tex_r0[46] ),
    .A1(\rbzero.tex_r0[45] ),
    .S(_04066_),
    .X(_04075_));
 sky130_fd_sc_hd__clkbuf_1 _10577_ (.A(_04075_),
    .X(_01515_));
 sky130_fd_sc_hd__mux2_1 _10578_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_04066_),
    .X(_04076_));
 sky130_fd_sc_hd__clkbuf_1 _10579_ (.A(_04076_),
    .X(_01514_));
 sky130_fd_sc_hd__clkbuf_4 _10580_ (.A(_04054_),
    .X(_04077_));
 sky130_fd_sc_hd__mux2_1 _10581_ (.A0(\rbzero.tex_r0[44] ),
    .A1(\rbzero.tex_r0[43] ),
    .S(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__clkbuf_1 _10582_ (.A(_04078_),
    .X(_01513_));
 sky130_fd_sc_hd__mux2_1 _10583_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_04077_),
    .X(_04079_));
 sky130_fd_sc_hd__clkbuf_1 _10584_ (.A(_04079_),
    .X(_01512_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(\rbzero.tex_r0[42] ),
    .A1(\rbzero.tex_r0[41] ),
    .S(_04077_),
    .X(_04080_));
 sky130_fd_sc_hd__clkbuf_1 _10586_ (.A(_04080_),
    .X(_01511_));
 sky130_fd_sc_hd__mux2_1 _10587_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_04077_),
    .X(_04081_));
 sky130_fd_sc_hd__clkbuf_1 _10588_ (.A(_04081_),
    .X(_01510_));
 sky130_fd_sc_hd__mux2_1 _10589_ (.A0(\rbzero.tex_r0[40] ),
    .A1(\rbzero.tex_r0[39] ),
    .S(_04077_),
    .X(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _10590_ (.A(_04082_),
    .X(_01509_));
 sky130_fd_sc_hd__mux2_1 _10591_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04077_),
    .X(_04083_));
 sky130_fd_sc_hd__clkbuf_1 _10592_ (.A(_04083_),
    .X(_01508_));
 sky130_fd_sc_hd__mux2_1 _10593_ (.A0(\rbzero.tex_r0[38] ),
    .A1(\rbzero.tex_r0[37] ),
    .S(_04077_),
    .X(_04084_));
 sky130_fd_sc_hd__clkbuf_1 _10594_ (.A(_04084_),
    .X(_01507_));
 sky130_fd_sc_hd__mux2_1 _10595_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_04077_),
    .X(_04085_));
 sky130_fd_sc_hd__clkbuf_1 _10596_ (.A(_04085_),
    .X(_01506_));
 sky130_fd_sc_hd__mux2_1 _10597_ (.A0(\rbzero.tex_r0[36] ),
    .A1(\rbzero.tex_r0[35] ),
    .S(_04077_),
    .X(_04086_));
 sky130_fd_sc_hd__clkbuf_1 _10598_ (.A(_04086_),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _10599_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_04077_),
    .X(_04087_));
 sky130_fd_sc_hd__clkbuf_1 _10600_ (.A(_04087_),
    .X(_01504_));
 sky130_fd_sc_hd__clkbuf_4 _10601_ (.A(_04054_),
    .X(_04088_));
 sky130_fd_sc_hd__mux2_1 _10602_ (.A0(\rbzero.tex_r0[34] ),
    .A1(\rbzero.tex_r0[33] ),
    .S(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__clkbuf_1 _10603_ (.A(_04089_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _10604_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_04088_),
    .X(_04090_));
 sky130_fd_sc_hd__clkbuf_1 _10605_ (.A(_04090_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _10606_ (.A0(\rbzero.tex_r0[32] ),
    .A1(\rbzero.tex_r0[31] ),
    .S(_04088_),
    .X(_04091_));
 sky130_fd_sc_hd__clkbuf_1 _10607_ (.A(_04091_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _10608_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_04088_),
    .X(_04092_));
 sky130_fd_sc_hd__clkbuf_1 _10609_ (.A(_04092_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _10610_ (.A0(\rbzero.tex_r0[30] ),
    .A1(\rbzero.tex_r0[29] ),
    .S(_04088_),
    .X(_04093_));
 sky130_fd_sc_hd__clkbuf_1 _10611_ (.A(_04093_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _10612_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_04088_),
    .X(_04094_));
 sky130_fd_sc_hd__clkbuf_1 _10613_ (.A(_04094_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _10614_ (.A0(\rbzero.tex_r0[28] ),
    .A1(\rbzero.tex_r0[27] ),
    .S(_04088_),
    .X(_04095_));
 sky130_fd_sc_hd__clkbuf_1 _10615_ (.A(_04095_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _10616_ (.A0(\rbzero.tex_r0[27] ),
    .A1(\rbzero.tex_r0[26] ),
    .S(_04088_),
    .X(_04096_));
 sky130_fd_sc_hd__clkbuf_1 _10617_ (.A(_04096_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(\rbzero.tex_r0[26] ),
    .A1(\rbzero.tex_r0[25] ),
    .S(_04088_),
    .X(_04097_));
 sky130_fd_sc_hd__clkbuf_1 _10619_ (.A(_04097_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_04088_),
    .X(_04098_));
 sky130_fd_sc_hd__clkbuf_1 _10621_ (.A(_04098_),
    .X(_01494_));
 sky130_fd_sc_hd__clkbuf_4 _10622_ (.A(_04054_),
    .X(_04099_));
 sky130_fd_sc_hd__mux2_1 _10623_ (.A0(\rbzero.tex_r0[24] ),
    .A1(\rbzero.tex_r0[23] ),
    .S(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_1 _10624_ (.A(_04100_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _10625_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_04099_),
    .X(_04101_));
 sky130_fd_sc_hd__clkbuf_1 _10626_ (.A(_04101_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _10627_ (.A0(\rbzero.tex_r0[22] ),
    .A1(\rbzero.tex_r0[21] ),
    .S(_04099_),
    .X(_04102_));
 sky130_fd_sc_hd__clkbuf_1 _10628_ (.A(_04102_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _10629_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_04099_),
    .X(_04103_));
 sky130_fd_sc_hd__clkbuf_1 _10630_ (.A(_04103_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _10631_ (.A0(\rbzero.tex_r0[20] ),
    .A1(\rbzero.tex_r0[19] ),
    .S(_04099_),
    .X(_04104_));
 sky130_fd_sc_hd__clkbuf_1 _10632_ (.A(_04104_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _10633_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_04099_),
    .X(_04105_));
 sky130_fd_sc_hd__clkbuf_1 _10634_ (.A(_04105_),
    .X(_01488_));
 sky130_fd_sc_hd__mux2_1 _10635_ (.A0(\rbzero.tex_r0[18] ),
    .A1(\rbzero.tex_r0[17] ),
    .S(_04099_),
    .X(_04106_));
 sky130_fd_sc_hd__clkbuf_1 _10636_ (.A(_04106_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _10637_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_04099_),
    .X(_04107_));
 sky130_fd_sc_hd__clkbuf_1 _10638_ (.A(_04107_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _10639_ (.A0(\rbzero.tex_r0[16] ),
    .A1(\rbzero.tex_r0[15] ),
    .S(_04099_),
    .X(_04108_));
 sky130_fd_sc_hd__clkbuf_1 _10640_ (.A(_04108_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _10641_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_04099_),
    .X(_04109_));
 sky130_fd_sc_hd__clkbuf_1 _10642_ (.A(_04109_),
    .X(_01484_));
 sky130_fd_sc_hd__clkbuf_4 _10643_ (.A(_04054_),
    .X(_04110_));
 sky130_fd_sc_hd__mux2_1 _10644_ (.A0(\rbzero.tex_r0[14] ),
    .A1(\rbzero.tex_r0[13] ),
    .S(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__clkbuf_1 _10645_ (.A(_04111_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _10646_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_04110_),
    .X(_04112_));
 sky130_fd_sc_hd__clkbuf_1 _10647_ (.A(_04112_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _10648_ (.A0(\rbzero.tex_r0[12] ),
    .A1(\rbzero.tex_r0[11] ),
    .S(_04110_),
    .X(_04113_));
 sky130_fd_sc_hd__clkbuf_1 _10649_ (.A(_04113_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_04110_),
    .X(_04114_));
 sky130_fd_sc_hd__clkbuf_1 _10651_ (.A(_04114_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _10652_ (.A0(\rbzero.tex_r0[10] ),
    .A1(\rbzero.tex_r0[9] ),
    .S(_04110_),
    .X(_04115_));
 sky130_fd_sc_hd__clkbuf_1 _10653_ (.A(_04115_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _10654_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_04110_),
    .X(_04116_));
 sky130_fd_sc_hd__clkbuf_1 _10655_ (.A(_04116_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _10656_ (.A0(\rbzero.tex_r0[8] ),
    .A1(\rbzero.tex_r0[7] ),
    .S(_04110_),
    .X(_04117_));
 sky130_fd_sc_hd__clkbuf_1 _10657_ (.A(_04117_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _10658_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_04110_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _10659_ (.A(_04118_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(\rbzero.tex_r0[6] ),
    .A1(\rbzero.tex_r0[5] ),
    .S(_04110_),
    .X(_04119_));
 sky130_fd_sc_hd__clkbuf_1 _10661_ (.A(_04119_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_04110_),
    .X(_04120_));
 sky130_fd_sc_hd__clkbuf_1 _10663_ (.A(_04120_),
    .X(_01474_));
 sky130_fd_sc_hd__clkbuf_4 _10664_ (.A(_04054_),
    .X(_04121_));
 sky130_fd_sc_hd__mux2_1 _10665_ (.A0(\rbzero.tex_r0[4] ),
    .A1(\rbzero.tex_r0[3] ),
    .S(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__clkbuf_1 _10666_ (.A(_04122_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _10667_ (.A0(\rbzero.tex_r0[3] ),
    .A1(\rbzero.tex_r0[2] ),
    .S(_04121_),
    .X(_04123_));
 sky130_fd_sc_hd__clkbuf_1 _10668_ (.A(_04123_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _10669_ (.A0(\rbzero.tex_r0[2] ),
    .A1(\rbzero.tex_r0[1] ),
    .S(_04121_),
    .X(_04124_));
 sky130_fd_sc_hd__clkbuf_1 _10670_ (.A(_04124_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _10671_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_04121_),
    .X(_04125_));
 sky130_fd_sc_hd__clkbuf_1 _10672_ (.A(_04125_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _10673_ (.A0(\rbzero.tex_g1[63] ),
    .A1(net50),
    .S(_04046_),
    .X(_04126_));
 sky130_fd_sc_hd__clkbuf_1 _10674_ (.A(_04126_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _10675_ (.A0(\rbzero.tex_g1[62] ),
    .A1(\rbzero.tex_g1[63] ),
    .S(_04046_),
    .X(_04127_));
 sky130_fd_sc_hd__clkbuf_1 _10676_ (.A(_04127_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _10677_ (.A0(\rbzero.tex_g1[61] ),
    .A1(\rbzero.tex_g1[62] ),
    .S(_04046_),
    .X(_04128_));
 sky130_fd_sc_hd__clkbuf_1 _10678_ (.A(_04128_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _10679_ (.A0(\rbzero.tex_g1[60] ),
    .A1(\rbzero.tex_g1[61] ),
    .S(_04046_),
    .X(_04129_));
 sky130_fd_sc_hd__clkbuf_1 _10680_ (.A(_04129_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _10681_ (.A0(\rbzero.tex_g1[59] ),
    .A1(\rbzero.tex_g1[60] ),
    .S(_04046_),
    .X(_04130_));
 sky130_fd_sc_hd__clkbuf_1 _10682_ (.A(_04130_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _10683_ (.A0(\rbzero.tex_g1[58] ),
    .A1(\rbzero.tex_g1[59] ),
    .S(_04046_),
    .X(_04131_));
 sky130_fd_sc_hd__clkbuf_1 _10684_ (.A(_04131_),
    .X(_01464_));
 sky130_fd_sc_hd__clkbuf_4 _10685_ (.A(_03979_),
    .X(_04132_));
 sky130_fd_sc_hd__mux2_1 _10686_ (.A0(\rbzero.tex_g1[57] ),
    .A1(\rbzero.tex_g1[58] ),
    .S(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_1 _10687_ (.A(_04133_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _10688_ (.A0(\rbzero.tex_g1[56] ),
    .A1(\rbzero.tex_g1[57] ),
    .S(_04132_),
    .X(_04134_));
 sky130_fd_sc_hd__clkbuf_1 _10689_ (.A(_04134_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _10690_ (.A0(\rbzero.tex_g1[55] ),
    .A1(\rbzero.tex_g1[56] ),
    .S(_04132_),
    .X(_04135_));
 sky130_fd_sc_hd__clkbuf_1 _10691_ (.A(_04135_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _10692_ (.A0(\rbzero.tex_g1[54] ),
    .A1(\rbzero.tex_g1[55] ),
    .S(_04132_),
    .X(_04136_));
 sky130_fd_sc_hd__clkbuf_1 _10693_ (.A(_04136_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _10694_ (.A0(\rbzero.tex_g1[53] ),
    .A1(\rbzero.tex_g1[54] ),
    .S(_04132_),
    .X(_04137_));
 sky130_fd_sc_hd__clkbuf_1 _10695_ (.A(_04137_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _10696_ (.A0(\rbzero.tex_g1[52] ),
    .A1(\rbzero.tex_g1[53] ),
    .S(_04132_),
    .X(_04138_));
 sky130_fd_sc_hd__clkbuf_1 _10697_ (.A(_04138_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(\rbzero.tex_g1[51] ),
    .A1(\rbzero.tex_g1[52] ),
    .S(_04132_),
    .X(_04139_));
 sky130_fd_sc_hd__clkbuf_1 _10699_ (.A(_04139_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _10700_ (.A0(\rbzero.tex_g1[50] ),
    .A1(\rbzero.tex_g1[51] ),
    .S(_04132_),
    .X(_04140_));
 sky130_fd_sc_hd__clkbuf_1 _10701_ (.A(_04140_),
    .X(_01456_));
 sky130_fd_sc_hd__mux2_1 _10702_ (.A0(\rbzero.tex_g1[49] ),
    .A1(\rbzero.tex_g1[50] ),
    .S(_04132_),
    .X(_04141_));
 sky130_fd_sc_hd__clkbuf_1 _10703_ (.A(_04141_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _10704_ (.A0(\rbzero.tex_g1[48] ),
    .A1(\rbzero.tex_g1[49] ),
    .S(_04132_),
    .X(_04142_));
 sky130_fd_sc_hd__clkbuf_1 _10705_ (.A(_04142_),
    .X(_01454_));
 sky130_fd_sc_hd__buf_4 _10706_ (.A(_03978_),
    .X(_04143_));
 sky130_fd_sc_hd__clkbuf_4 _10707_ (.A(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__mux2_1 _10708_ (.A0(\rbzero.tex_g1[47] ),
    .A1(\rbzero.tex_g1[48] ),
    .S(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__clkbuf_1 _10709_ (.A(_04145_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _10710_ (.A0(\rbzero.tex_g1[46] ),
    .A1(\rbzero.tex_g1[47] ),
    .S(_04144_),
    .X(_04146_));
 sky130_fd_sc_hd__clkbuf_1 _10711_ (.A(_04146_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _10712_ (.A0(\rbzero.tex_g1[45] ),
    .A1(\rbzero.tex_g1[46] ),
    .S(_04144_),
    .X(_04147_));
 sky130_fd_sc_hd__clkbuf_1 _10713_ (.A(_04147_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _10714_ (.A0(\rbzero.tex_g1[44] ),
    .A1(\rbzero.tex_g1[45] ),
    .S(_04144_),
    .X(_04148_));
 sky130_fd_sc_hd__clkbuf_1 _10715_ (.A(_04148_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(\rbzero.tex_g1[43] ),
    .A1(\rbzero.tex_g1[44] ),
    .S(_04144_),
    .X(_04149_));
 sky130_fd_sc_hd__clkbuf_1 _10717_ (.A(_04149_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _10718_ (.A0(\rbzero.tex_g1[42] ),
    .A1(\rbzero.tex_g1[43] ),
    .S(_04144_),
    .X(_04150_));
 sky130_fd_sc_hd__clkbuf_1 _10719_ (.A(_04150_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _10720_ (.A0(\rbzero.tex_g1[41] ),
    .A1(\rbzero.tex_g1[42] ),
    .S(_04144_),
    .X(_04151_));
 sky130_fd_sc_hd__clkbuf_1 _10721_ (.A(_04151_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _10722_ (.A0(\rbzero.tex_g1[40] ),
    .A1(\rbzero.tex_g1[41] ),
    .S(_04144_),
    .X(_04152_));
 sky130_fd_sc_hd__clkbuf_1 _10723_ (.A(_04152_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(\rbzero.tex_g1[39] ),
    .A1(\rbzero.tex_g1[40] ),
    .S(_04144_),
    .X(_04153_));
 sky130_fd_sc_hd__clkbuf_1 _10725_ (.A(_04153_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _10726_ (.A0(\rbzero.tex_g1[38] ),
    .A1(\rbzero.tex_g1[39] ),
    .S(_04144_),
    .X(_04154_));
 sky130_fd_sc_hd__clkbuf_1 _10727_ (.A(_04154_),
    .X(_01444_));
 sky130_fd_sc_hd__clkbuf_4 _10728_ (.A(_04143_),
    .X(_04155_));
 sky130_fd_sc_hd__mux2_1 _10729_ (.A0(\rbzero.tex_g1[37] ),
    .A1(\rbzero.tex_g1[38] ),
    .S(_04155_),
    .X(_04156_));
 sky130_fd_sc_hd__clkbuf_1 _10730_ (.A(_04156_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _10731_ (.A0(\rbzero.tex_g1[36] ),
    .A1(\rbzero.tex_g1[37] ),
    .S(_04155_),
    .X(_04157_));
 sky130_fd_sc_hd__clkbuf_1 _10732_ (.A(_04157_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _10733_ (.A0(\rbzero.tex_g1[35] ),
    .A1(\rbzero.tex_g1[36] ),
    .S(_04155_),
    .X(_04158_));
 sky130_fd_sc_hd__clkbuf_1 _10734_ (.A(_04158_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _10735_ (.A0(\rbzero.tex_g1[34] ),
    .A1(\rbzero.tex_g1[35] ),
    .S(_04155_),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_1 _10736_ (.A(_04159_),
    .X(_01440_));
 sky130_fd_sc_hd__mux2_1 _10737_ (.A0(\rbzero.tex_g1[33] ),
    .A1(\rbzero.tex_g1[34] ),
    .S(_04155_),
    .X(_04160_));
 sky130_fd_sc_hd__clkbuf_1 _10738_ (.A(_04160_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _10739_ (.A0(\rbzero.tex_g1[32] ),
    .A1(\rbzero.tex_g1[33] ),
    .S(_04155_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _10740_ (.A(_04161_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(\rbzero.tex_g1[31] ),
    .A1(\rbzero.tex_g1[32] ),
    .S(_04155_),
    .X(_04162_));
 sky130_fd_sc_hd__clkbuf_1 _10742_ (.A(_04162_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(\rbzero.tex_g1[30] ),
    .A1(\rbzero.tex_g1[31] ),
    .S(_04155_),
    .X(_04163_));
 sky130_fd_sc_hd__clkbuf_1 _10744_ (.A(_04163_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(\rbzero.tex_g1[29] ),
    .A1(\rbzero.tex_g1[30] ),
    .S(_04155_),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_1 _10746_ (.A(_04164_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _10747_ (.A0(\rbzero.tex_g1[28] ),
    .A1(\rbzero.tex_g1[29] ),
    .S(_04155_),
    .X(_04165_));
 sky130_fd_sc_hd__clkbuf_1 _10748_ (.A(_04165_),
    .X(_01434_));
 sky130_fd_sc_hd__clkbuf_4 _10749_ (.A(_04143_),
    .X(_04166_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(\rbzero.tex_g1[27] ),
    .A1(\rbzero.tex_g1[28] ),
    .S(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__clkbuf_1 _10751_ (.A(_04167_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(\rbzero.tex_g1[26] ),
    .A1(\rbzero.tex_g1[27] ),
    .S(_04166_),
    .X(_04168_));
 sky130_fd_sc_hd__clkbuf_1 _10753_ (.A(_04168_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(\rbzero.tex_g1[25] ),
    .A1(\rbzero.tex_g1[26] ),
    .S(_04166_),
    .X(_04169_));
 sky130_fd_sc_hd__clkbuf_1 _10755_ (.A(_04169_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(\rbzero.tex_g1[24] ),
    .A1(\rbzero.tex_g1[25] ),
    .S(_04166_),
    .X(_04170_));
 sky130_fd_sc_hd__clkbuf_1 _10757_ (.A(_04170_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(\rbzero.tex_g1[23] ),
    .A1(\rbzero.tex_g1[24] ),
    .S(_04166_),
    .X(_04171_));
 sky130_fd_sc_hd__clkbuf_1 _10759_ (.A(_04171_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(\rbzero.tex_g1[22] ),
    .A1(\rbzero.tex_g1[23] ),
    .S(_04166_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _10761_ (.A(_04172_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(\rbzero.tex_g1[21] ),
    .A1(\rbzero.tex_g1[22] ),
    .S(_04166_),
    .X(_04173_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(_04173_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(\rbzero.tex_g1[20] ),
    .A1(\rbzero.tex_g1[21] ),
    .S(_04166_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _10765_ (.A(_04174_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(\rbzero.tex_g1[19] ),
    .A1(\rbzero.tex_g1[20] ),
    .S(_04166_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _10767_ (.A(_04175_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(\rbzero.tex_g1[18] ),
    .A1(\rbzero.tex_g1[19] ),
    .S(_04166_),
    .X(_04176_));
 sky130_fd_sc_hd__clkbuf_1 _10769_ (.A(_04176_),
    .X(_01424_));
 sky130_fd_sc_hd__clkbuf_4 _10770_ (.A(_04143_),
    .X(_04177_));
 sky130_fd_sc_hd__mux2_1 _10771_ (.A0(\rbzero.tex_g1[17] ),
    .A1(\rbzero.tex_g1[18] ),
    .S(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _10772_ (.A(_04178_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _10773_ (.A0(\rbzero.tex_g1[16] ),
    .A1(\rbzero.tex_g1[17] ),
    .S(_04177_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _10774_ (.A(_04179_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _10775_ (.A0(\rbzero.tex_g1[15] ),
    .A1(\rbzero.tex_g1[16] ),
    .S(_04177_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _10776_ (.A(_04180_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(\rbzero.tex_g1[14] ),
    .A1(\rbzero.tex_g1[15] ),
    .S(_04177_),
    .X(_04181_));
 sky130_fd_sc_hd__clkbuf_1 _10778_ (.A(_04181_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(\rbzero.tex_g1[13] ),
    .A1(\rbzero.tex_g1[14] ),
    .S(_04177_),
    .X(_04182_));
 sky130_fd_sc_hd__clkbuf_1 _10780_ (.A(_04182_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(\rbzero.tex_g1[12] ),
    .A1(\rbzero.tex_g1[13] ),
    .S(_04177_),
    .X(_04183_));
 sky130_fd_sc_hd__clkbuf_1 _10782_ (.A(_04183_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(\rbzero.tex_g1[11] ),
    .A1(\rbzero.tex_g1[12] ),
    .S(_04177_),
    .X(_04184_));
 sky130_fd_sc_hd__clkbuf_1 _10784_ (.A(_04184_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(\rbzero.tex_g1[10] ),
    .A1(\rbzero.tex_g1[11] ),
    .S(_04177_),
    .X(_04185_));
 sky130_fd_sc_hd__clkbuf_1 _10786_ (.A(_04185_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(\rbzero.tex_g1[9] ),
    .A1(\rbzero.tex_g1[10] ),
    .S(_04177_),
    .X(_04186_));
 sky130_fd_sc_hd__clkbuf_1 _10788_ (.A(_04186_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(\rbzero.tex_g1[8] ),
    .A1(\rbzero.tex_g1[9] ),
    .S(_04177_),
    .X(_04187_));
 sky130_fd_sc_hd__clkbuf_1 _10790_ (.A(_04187_),
    .X(_01414_));
 sky130_fd_sc_hd__buf_4 _10791_ (.A(_04143_),
    .X(_04188_));
 sky130_fd_sc_hd__mux2_1 _10792_ (.A0(\rbzero.tex_g1[7] ),
    .A1(\rbzero.tex_g1[8] ),
    .S(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _10793_ (.A(_04189_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _10794_ (.A0(\rbzero.tex_g1[6] ),
    .A1(\rbzero.tex_g1[7] ),
    .S(_04188_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _10795_ (.A(_04190_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _10796_ (.A0(\rbzero.tex_g1[5] ),
    .A1(\rbzero.tex_g1[6] ),
    .S(_04188_),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _10797_ (.A(_04191_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _10798_ (.A0(\rbzero.tex_g1[4] ),
    .A1(\rbzero.tex_g1[5] ),
    .S(_04188_),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _10799_ (.A(_04192_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _10800_ (.A0(\rbzero.tex_g1[3] ),
    .A1(\rbzero.tex_g1[4] ),
    .S(_04188_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _10801_ (.A(_04193_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _10802_ (.A0(\rbzero.tex_g1[2] ),
    .A1(\rbzero.tex_g1[3] ),
    .S(_04188_),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_1 _10803_ (.A(_04194_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _10804_ (.A0(\rbzero.tex_g1[1] ),
    .A1(\rbzero.tex_g1[2] ),
    .S(_04188_),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _10805_ (.A(_04195_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _10806_ (.A0(\rbzero.tex_g1[0] ),
    .A1(\rbzero.tex_g1[1] ),
    .S(_04188_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _10807_ (.A(_04196_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(net50),
    .A1(\rbzero.tex_g0[63] ),
    .S(_04121_),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_1 _10809_ (.A(_04197_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(\rbzero.tex_g0[63] ),
    .A1(\rbzero.tex_g0[62] ),
    .S(_04121_),
    .X(_04198_));
 sky130_fd_sc_hd__clkbuf_1 _10811_ (.A(_04198_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _10812_ (.A0(\rbzero.tex_g0[62] ),
    .A1(\rbzero.tex_g0[61] ),
    .S(_04121_),
    .X(_04199_));
 sky130_fd_sc_hd__clkbuf_1 _10813_ (.A(_04199_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_04121_),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_1 _10815_ (.A(_04200_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(\rbzero.tex_g0[60] ),
    .A1(\rbzero.tex_g0[59] ),
    .S(_04121_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_1 _10817_ (.A(_04201_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_04121_),
    .X(_04202_));
 sky130_fd_sc_hd__clkbuf_1 _10819_ (.A(_04202_),
    .X(_01400_));
 sky130_fd_sc_hd__clkbuf_4 _10820_ (.A(_04054_),
    .X(_04203_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(\rbzero.tex_g0[58] ),
    .A1(\rbzero.tex_g0[57] ),
    .S(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__clkbuf_1 _10822_ (.A(_04204_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_04203_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_1 _10824_ (.A(_04205_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(\rbzero.tex_g0[56] ),
    .A1(\rbzero.tex_g0[55] ),
    .S(_04203_),
    .X(_04206_));
 sky130_fd_sc_hd__clkbuf_1 _10826_ (.A(_04206_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _10827_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_04203_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _10828_ (.A(_04207_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _10829_ (.A0(\rbzero.tex_g0[54] ),
    .A1(\rbzero.tex_g0[53] ),
    .S(_04203_),
    .X(_04208_));
 sky130_fd_sc_hd__clkbuf_1 _10830_ (.A(_04208_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_04203_),
    .X(_04209_));
 sky130_fd_sc_hd__clkbuf_1 _10832_ (.A(_04209_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(\rbzero.tex_g0[52] ),
    .A1(\rbzero.tex_g0[51] ),
    .S(_04203_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _10834_ (.A(_04210_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _10835_ (.A0(\rbzero.tex_g0[51] ),
    .A1(\rbzero.tex_g0[50] ),
    .S(_04203_),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _10836_ (.A(_04211_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _10837_ (.A0(\rbzero.tex_g0[50] ),
    .A1(\rbzero.tex_g0[49] ),
    .S(_04203_),
    .X(_04212_));
 sky130_fd_sc_hd__clkbuf_1 _10838_ (.A(_04212_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _10839_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_04203_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _10840_ (.A(_04213_),
    .X(_01390_));
 sky130_fd_sc_hd__buf_4 _10841_ (.A(_04053_),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_4 _10842_ (.A(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__mux2_1 _10843_ (.A0(\rbzero.tex_g0[48] ),
    .A1(\rbzero.tex_g0[47] ),
    .S(_04215_),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_1 _10844_ (.A(_04216_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _10845_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_04215_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _10846_ (.A(_04217_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _10847_ (.A0(\rbzero.tex_g0[46] ),
    .A1(\rbzero.tex_g0[45] ),
    .S(_04215_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _10848_ (.A(_04218_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_04215_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _10850_ (.A(_04219_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(\rbzero.tex_g0[44] ),
    .A1(\rbzero.tex_g0[43] ),
    .S(_04215_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_1 _10852_ (.A(_04220_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_04215_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _10854_ (.A(_04221_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(\rbzero.tex_g0[42] ),
    .A1(\rbzero.tex_g0[41] ),
    .S(_04215_),
    .X(_04222_));
 sky130_fd_sc_hd__clkbuf_1 _10856_ (.A(_04222_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_04215_),
    .X(_04223_));
 sky130_fd_sc_hd__clkbuf_1 _10858_ (.A(_04223_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _10859_ (.A0(\rbzero.tex_g0[40] ),
    .A1(\rbzero.tex_g0[39] ),
    .S(_04215_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(_04224_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_04215_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _10862_ (.A(_04225_),
    .X(_01380_));
 sky130_fd_sc_hd__clkbuf_4 _10863_ (.A(_04214_),
    .X(_04226_));
 sky130_fd_sc_hd__mux2_1 _10864_ (.A0(\rbzero.tex_g0[38] ),
    .A1(\rbzero.tex_g0[37] ),
    .S(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__clkbuf_1 _10865_ (.A(_04227_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _10866_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_04226_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_1 _10867_ (.A(_04228_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(\rbzero.tex_g0[36] ),
    .A1(\rbzero.tex_g0[35] ),
    .S(_04226_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _10869_ (.A(_04229_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _10870_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_04226_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _10871_ (.A(_04230_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _10872_ (.A0(\rbzero.tex_g0[34] ),
    .A1(\rbzero.tex_g0[33] ),
    .S(_04226_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _10873_ (.A(_04231_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _10874_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_04226_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _10875_ (.A(_04232_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _10876_ (.A0(\rbzero.tex_g0[32] ),
    .A1(\rbzero.tex_g0[31] ),
    .S(_04226_),
    .X(_04233_));
 sky130_fd_sc_hd__clkbuf_1 _10877_ (.A(_04233_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_04226_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_1 _10879_ (.A(_04234_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _10880_ (.A0(\rbzero.tex_g0[30] ),
    .A1(\rbzero.tex_g0[29] ),
    .S(_04226_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _10881_ (.A(_04235_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_04226_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_1 _10883_ (.A(_04236_),
    .X(_01370_));
 sky130_fd_sc_hd__clkbuf_4 _10884_ (.A(_04214_),
    .X(_04237_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(\rbzero.tex_g0[28] ),
    .A1(\rbzero.tex_g0[27] ),
    .S(_04237_),
    .X(_04238_));
 sky130_fd_sc_hd__clkbuf_1 _10886_ (.A(_04238_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _10887_ (.A0(\rbzero.tex_g0[27] ),
    .A1(\rbzero.tex_g0[26] ),
    .S(_04237_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _10888_ (.A(_04239_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(\rbzero.tex_g0[26] ),
    .A1(\rbzero.tex_g0[25] ),
    .S(_04237_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _10890_ (.A(_04240_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _10891_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_04237_),
    .X(_04241_));
 sky130_fd_sc_hd__clkbuf_1 _10892_ (.A(_04241_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(\rbzero.tex_g0[24] ),
    .A1(\rbzero.tex_g0[23] ),
    .S(_04237_),
    .X(_04242_));
 sky130_fd_sc_hd__clkbuf_1 _10894_ (.A(_04242_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _10895_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_04237_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_1 _10896_ (.A(_04243_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(\rbzero.tex_g0[22] ),
    .A1(\rbzero.tex_g0[21] ),
    .S(_04237_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _10898_ (.A(_04244_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_04237_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_1 _10900_ (.A(_04245_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(\rbzero.tex_g0[20] ),
    .A1(\rbzero.tex_g0[19] ),
    .S(_04237_),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _10902_ (.A(_04246_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_04237_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_1 _10904_ (.A(_04247_),
    .X(_01360_));
 sky130_fd_sc_hd__clkbuf_4 _10905_ (.A(_04214_),
    .X(_04248_));
 sky130_fd_sc_hd__mux2_1 _10906_ (.A0(\rbzero.tex_g0[18] ),
    .A1(\rbzero.tex_g0[17] ),
    .S(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_1 _10907_ (.A(_04249_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _10908_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_04248_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _10909_ (.A(_04250_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _10910_ (.A0(\rbzero.tex_g0[16] ),
    .A1(\rbzero.tex_g0[15] ),
    .S(_04248_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _10911_ (.A(_04251_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _10912_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_04248_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_1 _10913_ (.A(_04252_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _10914_ (.A0(\rbzero.tex_g0[14] ),
    .A1(\rbzero.tex_g0[13] ),
    .S(_04248_),
    .X(_04253_));
 sky130_fd_sc_hd__clkbuf_1 _10915_ (.A(_04253_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _10916_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_04248_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _10917_ (.A(_04254_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _10918_ (.A0(\rbzero.tex_g0[12] ),
    .A1(\rbzero.tex_g0[11] ),
    .S(_04248_),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_1 _10919_ (.A(_04255_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_04248_),
    .X(_04256_));
 sky130_fd_sc_hd__clkbuf_1 _10921_ (.A(_04256_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(\rbzero.tex_g0[10] ),
    .A1(\rbzero.tex_g0[9] ),
    .S(_04248_),
    .X(_04257_));
 sky130_fd_sc_hd__clkbuf_1 _10923_ (.A(_04257_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_04248_),
    .X(_04258_));
 sky130_fd_sc_hd__clkbuf_1 _10925_ (.A(_04258_),
    .X(_01350_));
 sky130_fd_sc_hd__buf_4 _10926_ (.A(_04214_),
    .X(_04259_));
 sky130_fd_sc_hd__mux2_1 _10927_ (.A0(\rbzero.tex_g0[8] ),
    .A1(\rbzero.tex_g0[7] ),
    .S(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__clkbuf_1 _10928_ (.A(_04260_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _10929_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_04259_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _10930_ (.A(_04261_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _10931_ (.A0(\rbzero.tex_g0[6] ),
    .A1(\rbzero.tex_g0[5] ),
    .S(_04259_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _10932_ (.A(_04262_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _10933_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_04259_),
    .X(_04263_));
 sky130_fd_sc_hd__clkbuf_1 _10934_ (.A(_04263_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _10935_ (.A0(\rbzero.tex_g0[4] ),
    .A1(\rbzero.tex_g0[3] ),
    .S(_04259_),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_1 _10936_ (.A(_04264_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _10937_ (.A0(\rbzero.tex_g0[3] ),
    .A1(\rbzero.tex_g0[2] ),
    .S(_04259_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _10938_ (.A(_04265_),
    .X(_01344_));
 sky130_fd_sc_hd__mux2_1 _10939_ (.A0(\rbzero.tex_g0[2] ),
    .A1(\rbzero.tex_g0[1] ),
    .S(_04259_),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_1 _10940_ (.A(_04266_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _10941_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_04259_),
    .X(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _10942_ (.A(_04267_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _10943_ (.A0(\rbzero.tex_b1[63] ),
    .A1(net51),
    .S(_04188_),
    .X(_04268_));
 sky130_fd_sc_hd__clkbuf_1 _10944_ (.A(_04268_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _10945_ (.A0(\rbzero.tex_b1[62] ),
    .A1(\rbzero.tex_b1[63] ),
    .S(_04188_),
    .X(_04269_));
 sky130_fd_sc_hd__clkbuf_1 _10946_ (.A(_04269_),
    .X(_01340_));
 sky130_fd_sc_hd__clkbuf_4 _10947_ (.A(_04143_),
    .X(_04270_));
 sky130_fd_sc_hd__mux2_1 _10948_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_04270_),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _10949_ (.A(_04271_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _10950_ (.A0(\rbzero.tex_b1[60] ),
    .A1(\rbzero.tex_b1[61] ),
    .S(_04270_),
    .X(_04272_));
 sky130_fd_sc_hd__clkbuf_1 _10951_ (.A(_04272_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _10952_ (.A0(\rbzero.tex_b1[59] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_04270_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_1 _10953_ (.A(_04273_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _10954_ (.A0(\rbzero.tex_b1[58] ),
    .A1(\rbzero.tex_b1[59] ),
    .S(_04270_),
    .X(_04274_));
 sky130_fd_sc_hd__clkbuf_1 _10955_ (.A(_04274_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _10956_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[58] ),
    .S(_04270_),
    .X(_04275_));
 sky130_fd_sc_hd__clkbuf_1 _10957_ (.A(_04275_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _10958_ (.A0(\rbzero.tex_b1[56] ),
    .A1(\rbzero.tex_b1[57] ),
    .S(_04270_),
    .X(_04276_));
 sky130_fd_sc_hd__clkbuf_1 _10959_ (.A(_04276_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_04270_),
    .X(_04277_));
 sky130_fd_sc_hd__clkbuf_1 _10961_ (.A(_04277_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _10962_ (.A0(\rbzero.tex_b1[54] ),
    .A1(\rbzero.tex_b1[55] ),
    .S(_04270_),
    .X(_04278_));
 sky130_fd_sc_hd__clkbuf_1 _10963_ (.A(_04278_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_04270_),
    .X(_04279_));
 sky130_fd_sc_hd__clkbuf_1 _10965_ (.A(_04279_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(\rbzero.tex_b1[52] ),
    .A1(\rbzero.tex_b1[53] ),
    .S(_04270_),
    .X(_04280_));
 sky130_fd_sc_hd__clkbuf_1 _10967_ (.A(_04280_),
    .X(_01330_));
 sky130_fd_sc_hd__clkbuf_4 _10968_ (.A(_04143_),
    .X(_04281_));
 sky130_fd_sc_hd__mux2_1 _10969_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_1 _10970_ (.A(_04282_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _10971_ (.A0(\rbzero.tex_b1[50] ),
    .A1(\rbzero.tex_b1[51] ),
    .S(_04281_),
    .X(_04283_));
 sky130_fd_sc_hd__clkbuf_1 _10972_ (.A(_04283_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _10973_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_04281_),
    .X(_04284_));
 sky130_fd_sc_hd__clkbuf_1 _10974_ (.A(_04284_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _10975_ (.A0(\rbzero.tex_b1[48] ),
    .A1(\rbzero.tex_b1[49] ),
    .S(_04281_),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_1 _10976_ (.A(_04285_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _10977_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_04281_),
    .X(_04286_));
 sky130_fd_sc_hd__clkbuf_1 _10978_ (.A(_04286_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _10979_ (.A0(\rbzero.tex_b1[46] ),
    .A1(\rbzero.tex_b1[47] ),
    .S(_04281_),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_1 _10980_ (.A(_04287_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _10981_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_04281_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_1 _10982_ (.A(_04288_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _10983_ (.A0(\rbzero.tex_b1[44] ),
    .A1(\rbzero.tex_b1[45] ),
    .S(_04281_),
    .X(_04289_));
 sky130_fd_sc_hd__clkbuf_1 _10984_ (.A(_04289_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _10985_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_04281_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _10986_ (.A(_04290_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _10987_ (.A0(\rbzero.tex_b1[42] ),
    .A1(\rbzero.tex_b1[43] ),
    .S(_04281_),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_1 _10988_ (.A(_04291_),
    .X(_01320_));
 sky130_fd_sc_hd__clkbuf_4 _10989_ (.A(_04143_),
    .X(_04292_));
 sky130_fd_sc_hd__mux2_1 _10990_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__clkbuf_1 _10991_ (.A(_04293_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _10992_ (.A0(\rbzero.tex_b1[40] ),
    .A1(\rbzero.tex_b1[41] ),
    .S(_04292_),
    .X(_04294_));
 sky130_fd_sc_hd__clkbuf_1 _10993_ (.A(_04294_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _10994_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_04292_),
    .X(_04295_));
 sky130_fd_sc_hd__clkbuf_1 _10995_ (.A(_04295_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _10996_ (.A0(\rbzero.tex_b1[38] ),
    .A1(\rbzero.tex_b1[39] ),
    .S(_04292_),
    .X(_04296_));
 sky130_fd_sc_hd__clkbuf_1 _10997_ (.A(_04296_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _10998_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_04292_),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_1 _10999_ (.A(_04297_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _11000_ (.A0(\rbzero.tex_b1[36] ),
    .A1(\rbzero.tex_b1[37] ),
    .S(_04292_),
    .X(_04298_));
 sky130_fd_sc_hd__clkbuf_1 _11001_ (.A(_04298_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _11002_ (.A0(\rbzero.tex_b1[35] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_04292_),
    .X(_04299_));
 sky130_fd_sc_hd__clkbuf_1 _11003_ (.A(_04299_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _11004_ (.A0(\rbzero.tex_b1[34] ),
    .A1(\rbzero.tex_b1[35] ),
    .S(_04292_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _11005_ (.A(_04300_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _11006_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[34] ),
    .S(_04292_),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_1 _11007_ (.A(_04301_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _11008_ (.A0(\rbzero.tex_b1[32] ),
    .A1(\rbzero.tex_b1[33] ),
    .S(_04292_),
    .X(_04302_));
 sky130_fd_sc_hd__clkbuf_1 _11009_ (.A(_04302_),
    .X(_01310_));
 sky130_fd_sc_hd__clkbuf_4 _11010_ (.A(_04143_),
    .X(_04303_));
 sky130_fd_sc_hd__mux2_1 _11011_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_04303_),
    .X(_04304_));
 sky130_fd_sc_hd__clkbuf_1 _11012_ (.A(_04304_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _11013_ (.A0(\rbzero.tex_b1[30] ),
    .A1(\rbzero.tex_b1[31] ),
    .S(_04303_),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_1 _11014_ (.A(_04305_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _11015_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_04303_),
    .X(_04306_));
 sky130_fd_sc_hd__clkbuf_1 _11016_ (.A(_04306_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _11017_ (.A0(\rbzero.tex_b1[28] ),
    .A1(\rbzero.tex_b1[29] ),
    .S(_04303_),
    .X(_04307_));
 sky130_fd_sc_hd__clkbuf_1 _11018_ (.A(_04307_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _11019_ (.A0(\rbzero.tex_b1[27] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_04303_),
    .X(_04308_));
 sky130_fd_sc_hd__clkbuf_1 _11020_ (.A(_04308_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(\rbzero.tex_b1[26] ),
    .A1(\rbzero.tex_b1[27] ),
    .S(_04303_),
    .X(_04309_));
 sky130_fd_sc_hd__clkbuf_1 _11022_ (.A(_04309_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _11023_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[26] ),
    .S(_04303_),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_1 _11024_ (.A(_04310_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _11025_ (.A0(\rbzero.tex_b1[24] ),
    .A1(\rbzero.tex_b1[25] ),
    .S(_04303_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_1 _11026_ (.A(_04311_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _11027_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_04303_),
    .X(_04312_));
 sky130_fd_sc_hd__clkbuf_1 _11028_ (.A(_04312_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _11029_ (.A0(\rbzero.tex_b1[22] ),
    .A1(\rbzero.tex_b1[23] ),
    .S(_04303_),
    .X(_04313_));
 sky130_fd_sc_hd__clkbuf_1 _11030_ (.A(_04313_),
    .X(_01300_));
 sky130_fd_sc_hd__clkbuf_4 _11031_ (.A(_04143_),
    .X(_04314_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_04314_),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_1 _11033_ (.A(_04315_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _11034_ (.A0(\rbzero.tex_b1[20] ),
    .A1(\rbzero.tex_b1[21] ),
    .S(_04314_),
    .X(_04316_));
 sky130_fd_sc_hd__clkbuf_1 _11035_ (.A(_04316_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _11036_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_04314_),
    .X(_04317_));
 sky130_fd_sc_hd__clkbuf_1 _11037_ (.A(_04317_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _11038_ (.A0(\rbzero.tex_b1[18] ),
    .A1(\rbzero.tex_b1[19] ),
    .S(_04314_),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_1 _11039_ (.A(_04318_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _11040_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_04314_),
    .X(_04319_));
 sky130_fd_sc_hd__clkbuf_1 _11041_ (.A(_04319_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _11042_ (.A0(\rbzero.tex_b1[16] ),
    .A1(\rbzero.tex_b1[17] ),
    .S(_04314_),
    .X(_04320_));
 sky130_fd_sc_hd__clkbuf_1 _11043_ (.A(_04320_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _11044_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_04314_),
    .X(_04321_));
 sky130_fd_sc_hd__clkbuf_1 _11045_ (.A(_04321_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _11046_ (.A0(\rbzero.tex_b1[14] ),
    .A1(\rbzero.tex_b1[15] ),
    .S(_04314_),
    .X(_04322_));
 sky130_fd_sc_hd__clkbuf_1 _11047_ (.A(_04322_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _11048_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_04314_),
    .X(_04323_));
 sky130_fd_sc_hd__clkbuf_1 _11049_ (.A(_04323_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _11050_ (.A0(\rbzero.tex_b1[12] ),
    .A1(\rbzero.tex_b1[13] ),
    .S(_04314_),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_1 _11051_ (.A(_04324_),
    .X(_01290_));
 sky130_fd_sc_hd__clkbuf_4 _11052_ (.A(_03978_),
    .X(_04325_));
 sky130_fd_sc_hd__mux2_1 _11053_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_04325_),
    .X(_04326_));
 sky130_fd_sc_hd__clkbuf_1 _11054_ (.A(_04326_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _11055_ (.A0(\rbzero.tex_b1[10] ),
    .A1(\rbzero.tex_b1[11] ),
    .S(_04325_),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_1 _11056_ (.A(_04327_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _11057_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_04325_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_1 _11058_ (.A(_04328_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _11059_ (.A0(\rbzero.tex_b1[8] ),
    .A1(\rbzero.tex_b1[9] ),
    .S(_04325_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _11060_ (.A(_04329_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _11061_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04325_),
    .X(_04330_));
 sky130_fd_sc_hd__clkbuf_1 _11062_ (.A(_04330_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _11063_ (.A0(\rbzero.tex_b1[6] ),
    .A1(\rbzero.tex_b1[7] ),
    .S(_04325_),
    .X(_04331_));
 sky130_fd_sc_hd__clkbuf_1 _11064_ (.A(_04331_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _11065_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_04325_),
    .X(_04332_));
 sky130_fd_sc_hd__clkbuf_1 _11066_ (.A(_04332_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _11067_ (.A0(\rbzero.tex_b1[4] ),
    .A1(\rbzero.tex_b1[5] ),
    .S(_04325_),
    .X(_04333_));
 sky130_fd_sc_hd__clkbuf_1 _11068_ (.A(_04333_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _11069_ (.A0(\rbzero.tex_b1[3] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_04325_),
    .X(_04334_));
 sky130_fd_sc_hd__clkbuf_1 _11070_ (.A(_04334_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _11071_ (.A0(\rbzero.tex_b1[2] ),
    .A1(\rbzero.tex_b1[3] ),
    .S(_04325_),
    .X(_04335_));
 sky130_fd_sc_hd__clkbuf_1 _11072_ (.A(_04335_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[2] ),
    .S(_03979_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _11074_ (.A(_04336_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _11075_ (.A0(\rbzero.tex_b1[0] ),
    .A1(\rbzero.tex_b1[1] ),
    .S(_03979_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_1 _11076_ (.A(_04337_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(net51),
    .A1(\rbzero.tex_b0[63] ),
    .S(_04259_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _11078_ (.A(_04338_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(\rbzero.tex_b0[63] ),
    .A1(\rbzero.tex_b0[62] ),
    .S(_04259_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _11080_ (.A(_04339_),
    .X(_01084_));
 sky130_fd_sc_hd__clkbuf_4 _11081_ (.A(_04214_),
    .X(_04340_));
 sky130_fd_sc_hd__mux2_1 _11082_ (.A0(\rbzero.tex_b0[62] ),
    .A1(\rbzero.tex_b0[61] ),
    .S(_04340_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_1 _11083_ (.A(_04341_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _11084_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_04340_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _11085_ (.A(_04342_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _11086_ (.A0(\rbzero.tex_b0[60] ),
    .A1(\rbzero.tex_b0[59] ),
    .S(_04340_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _11087_ (.A(_04343_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _11088_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_04340_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _11089_ (.A(_04344_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _11090_ (.A0(\rbzero.tex_b0[58] ),
    .A1(\rbzero.tex_b0[57] ),
    .S(_04340_),
    .X(_04345_));
 sky130_fd_sc_hd__clkbuf_1 _11091_ (.A(_04345_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _11092_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_04340_),
    .X(_04346_));
 sky130_fd_sc_hd__clkbuf_1 _11093_ (.A(_04346_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(\rbzero.tex_b0[56] ),
    .A1(\rbzero.tex_b0[55] ),
    .S(_04340_),
    .X(_04347_));
 sky130_fd_sc_hd__clkbuf_1 _11095_ (.A(_04347_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(\rbzero.tex_b0[55] ),
    .A1(\rbzero.tex_b0[54] ),
    .S(_04340_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _11097_ (.A(_04348_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(\rbzero.tex_b0[54] ),
    .A1(\rbzero.tex_b0[53] ),
    .S(_04340_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _11099_ (.A(_04349_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_04340_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_1 _11101_ (.A(_04350_),
    .X(_01074_));
 sky130_fd_sc_hd__clkbuf_4 _11102_ (.A(_04214_),
    .X(_04351_));
 sky130_fd_sc_hd__mux2_1 _11103_ (.A0(\rbzero.tex_b0[52] ),
    .A1(\rbzero.tex_b0[51] ),
    .S(_04351_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _11104_ (.A(_04352_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _11105_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_04351_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_1 _11106_ (.A(_04353_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _11107_ (.A0(\rbzero.tex_b0[50] ),
    .A1(\rbzero.tex_b0[49] ),
    .S(_04351_),
    .X(_04354_));
 sky130_fd_sc_hd__clkbuf_1 _11108_ (.A(_04354_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _11109_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_04351_),
    .X(_04355_));
 sky130_fd_sc_hd__clkbuf_1 _11110_ (.A(_04355_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _11111_ (.A0(\rbzero.tex_b0[48] ),
    .A1(\rbzero.tex_b0[47] ),
    .S(_04351_),
    .X(_04356_));
 sky130_fd_sc_hd__clkbuf_1 _11112_ (.A(_04356_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _11113_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_04351_),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _11114_ (.A(_04357_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(\rbzero.tex_b0[46] ),
    .A1(\rbzero.tex_b0[45] ),
    .S(_04351_),
    .X(_04358_));
 sky130_fd_sc_hd__clkbuf_1 _11116_ (.A(_04358_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_04351_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _11118_ (.A(_04359_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _11119_ (.A0(\rbzero.tex_b0[44] ),
    .A1(\rbzero.tex_b0[43] ),
    .S(_04351_),
    .X(_04360_));
 sky130_fd_sc_hd__clkbuf_1 _11120_ (.A(_04360_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _11121_ (.A0(\rbzero.tex_b0[43] ),
    .A1(\rbzero.tex_b0[42] ),
    .S(_04351_),
    .X(_04361_));
 sky130_fd_sc_hd__clkbuf_1 _11122_ (.A(_04361_),
    .X(_01064_));
 sky130_fd_sc_hd__clkbuf_4 _11123_ (.A(_04214_),
    .X(_04362_));
 sky130_fd_sc_hd__mux2_1 _11124_ (.A0(\rbzero.tex_b0[42] ),
    .A1(\rbzero.tex_b0[41] ),
    .S(_04362_),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _11125_ (.A(_04363_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _11126_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_04362_),
    .X(_04364_));
 sky130_fd_sc_hd__clkbuf_1 _11127_ (.A(_04364_),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _11128_ (.A0(\rbzero.tex_b0[40] ),
    .A1(\rbzero.tex_b0[39] ),
    .S(_04362_),
    .X(_04365_));
 sky130_fd_sc_hd__clkbuf_1 _11129_ (.A(_04365_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _11130_ (.A0(\rbzero.tex_b0[39] ),
    .A1(\rbzero.tex_b0[38] ),
    .S(_04362_),
    .X(_04366_));
 sky130_fd_sc_hd__clkbuf_1 _11131_ (.A(_04366_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _11132_ (.A0(\rbzero.tex_b0[38] ),
    .A1(\rbzero.tex_b0[37] ),
    .S(_04362_),
    .X(_04367_));
 sky130_fd_sc_hd__clkbuf_1 _11133_ (.A(_04367_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _11134_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_04362_),
    .X(_04368_));
 sky130_fd_sc_hd__clkbuf_1 _11135_ (.A(_04368_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _11136_ (.A0(\rbzero.tex_b0[36] ),
    .A1(\rbzero.tex_b0[35] ),
    .S(_04362_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_1 _11137_ (.A(_04369_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _11138_ (.A0(\rbzero.tex_b0[35] ),
    .A1(\rbzero.tex_b0[34] ),
    .S(_04362_),
    .X(_04370_));
 sky130_fd_sc_hd__clkbuf_1 _11139_ (.A(_04370_),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _11140_ (.A0(\rbzero.tex_b0[34] ),
    .A1(\rbzero.tex_b0[33] ),
    .S(_04362_),
    .X(_04371_));
 sky130_fd_sc_hd__clkbuf_1 _11141_ (.A(_04371_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _11142_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_04362_),
    .X(_04372_));
 sky130_fd_sc_hd__clkbuf_1 _11143_ (.A(_04372_),
    .X(_01054_));
 sky130_fd_sc_hd__clkbuf_4 _11144_ (.A(_04214_),
    .X(_04373_));
 sky130_fd_sc_hd__mux2_1 _11145_ (.A0(\rbzero.tex_b0[32] ),
    .A1(\rbzero.tex_b0[31] ),
    .S(_04373_),
    .X(_04374_));
 sky130_fd_sc_hd__clkbuf_1 _11146_ (.A(_04374_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _11147_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_04373_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_1 _11148_ (.A(_04375_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _11149_ (.A0(\rbzero.tex_b0[30] ),
    .A1(\rbzero.tex_b0[29] ),
    .S(_04373_),
    .X(_04376_));
 sky130_fd_sc_hd__clkbuf_1 _11150_ (.A(_04376_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _11151_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_04373_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_1 _11152_ (.A(_04377_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _11153_ (.A0(\rbzero.tex_b0[28] ),
    .A1(\rbzero.tex_b0[27] ),
    .S(_04373_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_1 _11154_ (.A(_04378_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _11155_ (.A0(\rbzero.tex_b0[27] ),
    .A1(\rbzero.tex_b0[26] ),
    .S(_04373_),
    .X(_04379_));
 sky130_fd_sc_hd__clkbuf_1 _11156_ (.A(_04379_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _11157_ (.A0(\rbzero.tex_b0[26] ),
    .A1(\rbzero.tex_b0[25] ),
    .S(_04373_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_1 _11158_ (.A(_04380_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _11159_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_04373_),
    .X(_04381_));
 sky130_fd_sc_hd__clkbuf_1 _11160_ (.A(_04381_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _11161_ (.A0(\rbzero.tex_b0[24] ),
    .A1(\rbzero.tex_b0[23] ),
    .S(_04373_),
    .X(_04382_));
 sky130_fd_sc_hd__clkbuf_1 _11162_ (.A(_04382_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _11163_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_04373_),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_1 _11164_ (.A(_04383_),
    .X(_01044_));
 sky130_fd_sc_hd__clkbuf_4 _11165_ (.A(_04214_),
    .X(_04384_));
 sky130_fd_sc_hd__mux2_1 _11166_ (.A0(\rbzero.tex_b0[22] ),
    .A1(\rbzero.tex_b0[21] ),
    .S(_04384_),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_1 _11167_ (.A(_04385_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _11168_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_04384_),
    .X(_04386_));
 sky130_fd_sc_hd__clkbuf_1 _11169_ (.A(_04386_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _11170_ (.A0(\rbzero.tex_b0[20] ),
    .A1(\rbzero.tex_b0[19] ),
    .S(_04384_),
    .X(_04387_));
 sky130_fd_sc_hd__clkbuf_1 _11171_ (.A(_04387_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _11172_ (.A0(\rbzero.tex_b0[19] ),
    .A1(\rbzero.tex_b0[18] ),
    .S(_04384_),
    .X(_04388_));
 sky130_fd_sc_hd__clkbuf_1 _11173_ (.A(_04388_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _11174_ (.A0(\rbzero.tex_b0[18] ),
    .A1(\rbzero.tex_b0[17] ),
    .S(_04384_),
    .X(_04389_));
 sky130_fd_sc_hd__clkbuf_1 _11175_ (.A(_04389_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _11176_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_04384_),
    .X(_04390_));
 sky130_fd_sc_hd__clkbuf_1 _11177_ (.A(_04390_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _11178_ (.A0(\rbzero.tex_b0[16] ),
    .A1(\rbzero.tex_b0[15] ),
    .S(_04384_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _11179_ (.A(_04391_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _11180_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_04384_),
    .X(_04392_));
 sky130_fd_sc_hd__clkbuf_1 _11181_ (.A(_04392_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _11182_ (.A0(\rbzero.tex_b0[14] ),
    .A1(\rbzero.tex_b0[13] ),
    .S(_04384_),
    .X(_04393_));
 sky130_fd_sc_hd__clkbuf_1 _11183_ (.A(_04393_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _11184_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_04384_),
    .X(_04394_));
 sky130_fd_sc_hd__clkbuf_1 _11185_ (.A(_04394_),
    .X(_01034_));
 sky130_fd_sc_hd__clkbuf_4 _11186_ (.A(_04053_),
    .X(_04395_));
 sky130_fd_sc_hd__mux2_1 _11187_ (.A0(\rbzero.tex_b0[12] ),
    .A1(\rbzero.tex_b0[11] ),
    .S(_04395_),
    .X(_04396_));
 sky130_fd_sc_hd__clkbuf_1 _11188_ (.A(_04396_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _11189_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_04395_),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_1 _11190_ (.A(_04397_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _11191_ (.A0(\rbzero.tex_b0[10] ),
    .A1(\rbzero.tex_b0[9] ),
    .S(_04395_),
    .X(_04398_));
 sky130_fd_sc_hd__clkbuf_1 _11192_ (.A(_04398_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _11193_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_04395_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_1 _11194_ (.A(_04399_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _11195_ (.A0(\rbzero.tex_b0[8] ),
    .A1(\rbzero.tex_b0[7] ),
    .S(_04395_),
    .X(_04400_));
 sky130_fd_sc_hd__clkbuf_1 _11196_ (.A(_04400_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _11197_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_04395_),
    .X(_04401_));
 sky130_fd_sc_hd__clkbuf_1 _11198_ (.A(_04401_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _11199_ (.A0(\rbzero.tex_b0[6] ),
    .A1(\rbzero.tex_b0[5] ),
    .S(_04395_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _11200_ (.A(_04402_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _11201_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_04395_),
    .X(_04403_));
 sky130_fd_sc_hd__clkbuf_1 _11202_ (.A(_04403_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _11203_ (.A0(\rbzero.tex_b0[4] ),
    .A1(\rbzero.tex_b0[3] ),
    .S(_04395_),
    .X(_04404_));
 sky130_fd_sc_hd__clkbuf_1 _11204_ (.A(_04404_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _11205_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_04395_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _11206_ (.A(_04405_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(\rbzero.tex_b0[2] ),
    .A1(\rbzero.tex_b0[1] ),
    .S(_04054_),
    .X(_04406_));
 sky130_fd_sc_hd__clkbuf_1 _11208_ (.A(_04406_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _11209_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_04054_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_1 _11210_ (.A(_04407_),
    .X(_01022_));
 sky130_fd_sc_hd__buf_6 _11211_ (.A(_04052_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_8 _11212_ (.A(_04408_),
    .X(_04409_));
 sky130_fd_sc_hd__buf_8 _11213_ (.A(_04409_),
    .X(net63));
 sky130_fd_sc_hd__inv_2 _11214_ (.A(\gpout0.hpos[6] ),
    .Y(_04410_));
 sky130_fd_sc_hd__buf_4 _11215_ (.A(\gpout0.hpos[5] ),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_4 _11216_ (.A(\gpout0.hpos[3] ),
    .X(_04412_));
 sky130_fd_sc_hd__inv_2 _11217_ (.A(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__inv_4 _11218_ (.A(\gpout0.hpos[4] ),
    .Y(_04414_));
 sky130_fd_sc_hd__nor2_2 _11219_ (.A(_04413_),
    .B(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__nor2_1 _11220_ (.A(_04411_),
    .B(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__o21ai_2 _11221_ (.A1(_04410_),
    .A2(_04416_),
    .B1(_04051_),
    .Y(_04417_));
 sky130_fd_sc_hd__buf_4 _11222_ (.A(\gpout0.hpos[6] ),
    .X(_04418_));
 sky130_fd_sc_hd__clkbuf_4 _11223_ (.A(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__buf_4 _11224_ (.A(\gpout0.hpos[9] ),
    .X(_04420_));
 sky130_fd_sc_hd__clkinv_2 _11225_ (.A(\gpout0.hpos[5] ),
    .Y(_04421_));
 sky130_fd_sc_hd__nand2_1 _11226_ (.A(_04412_),
    .B(\gpout0.hpos[4] ),
    .Y(_04422_));
 sky130_fd_sc_hd__nor2_1 _11227_ (.A(_04421_),
    .B(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hd__nor2_2 _11228_ (.A(_04416_),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__and4_1 _11229_ (.A(_04051_),
    .B(_04419_),
    .C(_04420_),
    .D(_04424_),
    .X(_04425_));
 sky130_fd_sc_hd__a21boi_2 _11230_ (.A1(_03975_),
    .A2(_04417_),
    .B1_N(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__inv_4 _11231_ (.A(_04426_),
    .Y(net71));
 sky130_fd_sc_hd__buf_2 _11232_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_04427_));
 sky130_fd_sc_hd__buf_2 _11233_ (.A(_04427_),
    .X(_04428_));
 sky130_fd_sc_hd__buf_4 _11234_ (.A(\rbzero.trace_state[2] ),
    .X(_04429_));
 sky130_fd_sc_hd__or2_2 _11235_ (.A(\rbzero.trace_state[1] ),
    .B(\rbzero.trace_state[0] ),
    .X(_04430_));
 sky130_fd_sc_hd__inv_2 _11236_ (.A(\rbzero.vga_sync.vsync ),
    .Y(_04431_));
 sky130_fd_sc_hd__nand2_4 _11237_ (.A(_04431_),
    .B(_03974_),
    .Y(_04432_));
 sky130_fd_sc_hd__inv_4 _11238_ (.A(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__buf_4 _11239_ (.A(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__o31a_1 _11240_ (.A1(\rbzero.trace_state[3] ),
    .A2(_04429_),
    .A3(_04430_),
    .B1(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__buf_4 _11241_ (.A(\rbzero.trace_state[1] ),
    .X(_04436_));
 sky130_fd_sc_hd__buf_2 _11242_ (.A(\rbzero.trace_state[0] ),
    .X(_04437_));
 sky130_fd_sc_hd__nor2_1 _11243_ (.A(\rbzero.trace_state[3] ),
    .B(_04429_),
    .Y(_04438_));
 sky130_fd_sc_hd__and3_1 _11244_ (.A(_04436_),
    .B(_04437_),
    .C(_04438_),
    .X(_04439_));
 sky130_fd_sc_hd__and4bb_1 _11245_ (.A_N(_04429_),
    .B_N(_04436_),
    .C(_04437_),
    .D(\rbzero.trace_state[3] ),
    .X(_04440_));
 sky130_fd_sc_hd__nor2_1 _11246_ (.A(_04439_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__clkbuf_8 _11247_ (.A(_04434_),
    .X(_04442_));
 sky130_fd_sc_hd__a32o_1 _11248_ (.A1(_04428_),
    .A2(_04435_),
    .A3(_04441_),
    .B1(_04439_),
    .B2(_04442_),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_2 _11249_ (.A(_03977_),
    .B(_04417_),
    .Y(net70));
 sky130_fd_sc_hd__clkbuf_4 _11250_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_04443_));
 sky130_fd_sc_hd__buf_2 _11251_ (.A(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__a21bo_1 _11252_ (.A1(_04444_),
    .A2(_04441_),
    .B1_N(_04435_),
    .X(_00000_));
 sky130_fd_sc_hd__inv_2 _11253_ (.A(\gpout0.hpos[2] ),
    .Y(_04445_));
 sky130_fd_sc_hd__buf_4 _11254_ (.A(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__or2_1 _11255_ (.A(\gpout0.hpos[1] ),
    .B(\gpout0.hpos[0] ),
    .X(_04447_));
 sky130_fd_sc_hd__nand2_2 _11256_ (.A(\gpout0.hpos[1] ),
    .B(\gpout0.hpos[0] ),
    .Y(_04448_));
 sky130_fd_sc_hd__inv_4 _11257_ (.A(\gpout0.hpos[1] ),
    .Y(_04449_));
 sky130_fd_sc_hd__a21oi_1 _11258_ (.A1(_04449_),
    .A2(_03971_),
    .B1(_04446_),
    .Y(_04450_));
 sky130_fd_sc_hd__a31o_1 _11259_ (.A1(_04446_),
    .A2(_04447_),
    .A3(_04448_),
    .B1(_04450_),
    .X(_04451_));
 sky130_fd_sc_hd__buf_4 _11260_ (.A(\gpout0.hpos[2] ),
    .X(_04452_));
 sky130_fd_sc_hd__inv_2 _11261_ (.A(_03969_),
    .Y(_04453_));
 sky130_fd_sc_hd__buf_4 _11262_ (.A(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__and2_1 _11263_ (.A(\rbzero.wall_hot[1] ),
    .B(\rbzero.wall_hot[0] ),
    .X(_04455_));
 sky130_fd_sc_hd__clkbuf_4 _11264_ (.A(_04455_),
    .X(_04456_));
 sky130_fd_sc_hd__nor2_4 _11265_ (.A(\rbzero.wall_hot[1] ),
    .B(\rbzero.wall_hot[0] ),
    .Y(_04457_));
 sky130_fd_sc_hd__a22o_1 _11266_ (.A1(\rbzero.spi_registers.texadd2[14] ),
    .A2(_04456_),
    .B1(_04457_),
    .B2(\rbzero.spi_registers.texadd3[14] ),
    .X(_04458_));
 sky130_fd_sc_hd__inv_2 _11267_ (.A(\rbzero.wall_hot[1] ),
    .Y(_04459_));
 sky130_fd_sc_hd__nor2_2 _11268_ (.A(_04459_),
    .B(\rbzero.wall_hot[0] ),
    .Y(_04460_));
 sky130_fd_sc_hd__clkbuf_4 _11269_ (.A(_04460_),
    .X(_04461_));
 sky130_fd_sc_hd__a22o_1 _11270_ (.A1(\rbzero.spi_registers.texadd3[13] ),
    .A2(_04457_),
    .B1(_04461_),
    .B2(\rbzero.spi_registers.texadd1[13] ),
    .X(_04462_));
 sky130_fd_sc_hd__buf_2 _11271_ (.A(\rbzero.side_hot ),
    .X(_04463_));
 sky130_fd_sc_hd__buf_4 _11272_ (.A(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__clkbuf_4 _11273_ (.A(_04459_),
    .X(_04465_));
 sky130_fd_sc_hd__nand2_1 _11274_ (.A(_04465_),
    .B(\rbzero.wall_hot[0] ),
    .Y(_04466_));
 sky130_fd_sc_hd__clkbuf_4 _11275_ (.A(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__and2_1 _11276_ (.A(\rbzero.spi_registers.texadd1[12] ),
    .B(_04461_),
    .X(_04468_));
 sky130_fd_sc_hd__and2_1 _11277_ (.A(_04459_),
    .B(\rbzero.wall_hot[0] ),
    .X(_04469_));
 sky130_fd_sc_hd__clkbuf_4 _11278_ (.A(_04469_),
    .X(_04470_));
 sky130_fd_sc_hd__a221o_1 _11279_ (.A1(\rbzero.spi_registers.texadd3[12] ),
    .A2(_04465_),
    .B1(_04456_),
    .B2(\rbzero.spi_registers.texadd2[12] ),
    .C1(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__o22a_1 _11280_ (.A1(\rbzero.spi_registers.texadd0[12] ),
    .A2(_04467_),
    .B1(_04468_),
    .B2(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__and2_1 _11281_ (.A(_04464_),
    .B(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__and2_1 _11282_ (.A(\rbzero.spi_registers.texadd1[11] ),
    .B(_04461_),
    .X(_04474_));
 sky130_fd_sc_hd__a221o_1 _11283_ (.A1(\rbzero.spi_registers.texadd3[11] ),
    .A2(_04465_),
    .B1(_04456_),
    .B2(\rbzero.spi_registers.texadd2[11] ),
    .C1(_04470_),
    .X(_04475_));
 sky130_fd_sc_hd__o22a_1 _11284_ (.A1(\rbzero.spi_registers.texadd0[11] ),
    .A2(_04467_),
    .B1(_04474_),
    .B2(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__nand2_1 _11285_ (.A(\rbzero.texu_hot[5] ),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__and2_1 _11286_ (.A(\rbzero.spi_registers.texadd1[10] ),
    .B(_04460_),
    .X(_04478_));
 sky130_fd_sc_hd__a221o_1 _11287_ (.A1(\rbzero.spi_registers.texadd3[10] ),
    .A2(_04465_),
    .B1(_04456_),
    .B2(\rbzero.spi_registers.texadd2[10] ),
    .C1(_04470_),
    .X(_04479_));
 sky130_fd_sc_hd__o22a_1 _11288_ (.A1(\rbzero.spi_registers.texadd0[10] ),
    .A2(_04467_),
    .B1(_04478_),
    .B2(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__nand2_1 _11289_ (.A(\rbzero.texu_hot[4] ),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__and2_1 _11290_ (.A(\rbzero.spi_registers.texadd1[9] ),
    .B(_04460_),
    .X(_04482_));
 sky130_fd_sc_hd__a221o_1 _11291_ (.A1(\rbzero.spi_registers.texadd3[9] ),
    .A2(_04465_),
    .B1(_04456_),
    .B2(\rbzero.spi_registers.texadd2[9] ),
    .C1(_04470_),
    .X(_04483_));
 sky130_fd_sc_hd__o22a_1 _11292_ (.A1(\rbzero.spi_registers.texadd0[9] ),
    .A2(_04467_),
    .B1(_04482_),
    .B2(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__nand2_1 _11293_ (.A(\rbzero.texu_hot[3] ),
    .B(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__a22o_1 _11294_ (.A1(\rbzero.spi_registers.texadd3[8] ),
    .A2(_04465_),
    .B1(_04455_),
    .B2(\rbzero.spi_registers.texadd2[8] ),
    .X(_04486_));
 sky130_fd_sc_hd__a211o_1 _11295_ (.A1(\rbzero.spi_registers.texadd1[8] ),
    .A2(_04460_),
    .B1(_04470_),
    .C1(_04486_),
    .X(_04487_));
 sky130_fd_sc_hd__o21a_1 _11296_ (.A1(\rbzero.spi_registers.texadd0[8] ),
    .A2(_04466_),
    .B1(_04487_),
    .X(_04488_));
 sky130_fd_sc_hd__xnor2_1 _11297_ (.A(\rbzero.texu_hot[2] ),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__and2_1 _11298_ (.A(\rbzero.spi_registers.texadd1[7] ),
    .B(_04460_),
    .X(_04490_));
 sky130_fd_sc_hd__a221o_1 _11299_ (.A1(\rbzero.spi_registers.texadd3[7] ),
    .A2(_04465_),
    .B1(_04455_),
    .B2(\rbzero.spi_registers.texadd2[7] ),
    .C1(_04469_),
    .X(_04491_));
 sky130_fd_sc_hd__o22a_1 _11300_ (.A1(\rbzero.spi_registers.texadd0[7] ),
    .A2(_04466_),
    .B1(_04490_),
    .B2(_04491_),
    .X(_04492_));
 sky130_fd_sc_hd__a22o_1 _11301_ (.A1(\rbzero.spi_registers.texadd3[6] ),
    .A2(_04465_),
    .B1(_04455_),
    .B2(\rbzero.spi_registers.texadd2[6] ),
    .X(_04493_));
 sky130_fd_sc_hd__a211o_1 _11302_ (.A1(\rbzero.spi_registers.texadd1[6] ),
    .A2(_04460_),
    .B1(_04469_),
    .C1(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__or2_1 _11303_ (.A(\rbzero.spi_registers.texadd0[6] ),
    .B(_04466_),
    .X(_04495_));
 sky130_fd_sc_hd__nand3_1 _11304_ (.A(\rbzero.texu_hot[0] ),
    .B(_04494_),
    .C(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__xnor2_1 _11305_ (.A(\rbzero.texu_hot[1] ),
    .B(_04492_),
    .Y(_04497_));
 sky130_fd_sc_hd__nor2_1 _11306_ (.A(_04496_),
    .B(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hd__a21o_1 _11307_ (.A1(\rbzero.texu_hot[1] ),
    .A2(_04492_),
    .B1(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__and2b_1 _11308_ (.A_N(_04489_),
    .B(_04499_),
    .X(_04500_));
 sky130_fd_sc_hd__a21oi_1 _11309_ (.A1(\rbzero.texu_hot[2] ),
    .A2(_04488_),
    .B1(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__or2_1 _11310_ (.A(\rbzero.texu_hot[3] ),
    .B(_04484_),
    .X(_04502_));
 sky130_fd_sc_hd__nand2_1 _11311_ (.A(_04485_),
    .B(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__or2_1 _11312_ (.A(_04501_),
    .B(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__or2_1 _11313_ (.A(\rbzero.texu_hot[4] ),
    .B(_04480_),
    .X(_04505_));
 sky130_fd_sc_hd__nand2_1 _11314_ (.A(_04481_),
    .B(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__a21o_1 _11315_ (.A1(_04485_),
    .A2(_04504_),
    .B1(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__or2_1 _11316_ (.A(\rbzero.texu_hot[5] ),
    .B(_04476_),
    .X(_04508_));
 sky130_fd_sc_hd__nand2_1 _11317_ (.A(_04477_),
    .B(_04508_),
    .Y(_04509_));
 sky130_fd_sc_hd__a21o_1 _11318_ (.A1(_04481_),
    .A2(_04507_),
    .B1(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__nor2_1 _11319_ (.A(_04464_),
    .B(_04472_),
    .Y(_04511_));
 sky130_fd_sc_hd__or2_1 _11320_ (.A(_04473_),
    .B(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__a21oi_1 _11321_ (.A1(_04477_),
    .A2(_04510_),
    .B1(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__inv_2 _11322_ (.A(\rbzero.spi_registers.texadd2[13] ),
    .Y(_04514_));
 sky130_fd_sc_hd__a21oi_1 _11323_ (.A1(_04514_),
    .A2(_04456_),
    .B1(_04462_),
    .Y(_04515_));
 sky130_fd_sc_hd__o21a_1 _11324_ (.A1(\rbzero.spi_registers.texadd0[13] ),
    .A2(_04467_),
    .B1(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__o21a_1 _11325_ (.A1(_04473_),
    .A2(_04513_),
    .B1(_04516_),
    .X(_04517_));
 sky130_fd_sc_hd__or2_1 _11326_ (.A(\rbzero.spi_registers.texadd0[14] ),
    .B(_04467_),
    .X(_04518_));
 sky130_fd_sc_hd__inv_2 _11327_ (.A(\rbzero.spi_registers.texadd1[14] ),
    .Y(_04519_));
 sky130_fd_sc_hd__a21oi_1 _11328_ (.A1(_04519_),
    .A2(_04461_),
    .B1(_04458_),
    .Y(_04520_));
 sky130_fd_sc_hd__o211a_1 _11329_ (.A1(_04462_),
    .A2(_04517_),
    .B1(_04518_),
    .C1(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__a22o_1 _11330_ (.A1(\rbzero.spi_registers.texadd3[15] ),
    .A2(_04465_),
    .B1(_04456_),
    .B2(\rbzero.spi_registers.texadd2[15] ),
    .X(_04522_));
 sky130_fd_sc_hd__a211o_1 _11331_ (.A1(\rbzero.spi_registers.texadd1[15] ),
    .A2(_04461_),
    .B1(_04470_),
    .C1(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__o21a_1 _11332_ (.A1(\rbzero.spi_registers.texadd0[15] ),
    .A2(_04467_),
    .B1(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__o21ai_1 _11333_ (.A1(_04458_),
    .A2(_04521_),
    .B1(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__buf_4 _11334_ (.A(_04465_),
    .X(_04526_));
 sky130_fd_sc_hd__a22o_1 _11335_ (.A1(\rbzero.spi_registers.texadd3[16] ),
    .A2(_04526_),
    .B1(_04456_),
    .B2(\rbzero.spi_registers.texadd2[16] ),
    .X(_04527_));
 sky130_fd_sc_hd__a211o_1 _11336_ (.A1(\rbzero.spi_registers.texadd1[16] ),
    .A2(_04461_),
    .B1(_04470_),
    .C1(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__o21ai_1 _11337_ (.A1(\rbzero.spi_registers.texadd0[16] ),
    .A2(_04467_),
    .B1(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__nor2_1 _11338_ (.A(_04525_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__a22o_1 _11339_ (.A1(\rbzero.spi_registers.texadd3[17] ),
    .A2(_04526_),
    .B1(_04456_),
    .B2(\rbzero.spi_registers.texadd2[17] ),
    .X(_04531_));
 sky130_fd_sc_hd__a211o_1 _11340_ (.A1(\rbzero.spi_registers.texadd1[17] ),
    .A2(_04461_),
    .B1(_04470_),
    .C1(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__o21a_1 _11341_ (.A1(\rbzero.spi_registers.texadd0[17] ),
    .A2(_04467_),
    .B1(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__and2_1 _11342_ (.A(_04530_),
    .B(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__clkbuf_4 _11343_ (.A(_04467_),
    .X(_04535_));
 sky130_fd_sc_hd__clkbuf_4 _11344_ (.A(_04470_),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_4 _11345_ (.A(_04456_),
    .X(_04537_));
 sky130_fd_sc_hd__a22o_1 _11346_ (.A1(\rbzero.spi_registers.texadd3[18] ),
    .A2(_04526_),
    .B1(_04537_),
    .B2(\rbzero.spi_registers.texadd2[18] ),
    .X(_04538_));
 sky130_fd_sc_hd__a211o_1 _11347_ (.A1(\rbzero.spi_registers.texadd1[18] ),
    .A2(_04461_),
    .B1(_04536_),
    .C1(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__o21a_1 _11348_ (.A1(\rbzero.spi_registers.texadd0[18] ),
    .A2(_04535_),
    .B1(_04539_),
    .X(_04540_));
 sky130_fd_sc_hd__a22o_1 _11349_ (.A1(\rbzero.spi_registers.texadd3[19] ),
    .A2(_04526_),
    .B1(_04537_),
    .B2(\rbzero.spi_registers.texadd2[19] ),
    .X(_04541_));
 sky130_fd_sc_hd__a211o_1 _11350_ (.A1(\rbzero.spi_registers.texadd1[19] ),
    .A2(_04461_),
    .B1(_04470_),
    .C1(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__o21a_1 _11351_ (.A1(\rbzero.spi_registers.texadd0[19] ),
    .A2(_04535_),
    .B1(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__and3_1 _11352_ (.A(_04534_),
    .B(_04540_),
    .C(_04543_),
    .X(_04544_));
 sky130_fd_sc_hd__clkbuf_4 _11353_ (.A(_04461_),
    .X(_04545_));
 sky130_fd_sc_hd__a22o_1 _11354_ (.A1(\rbzero.spi_registers.texadd3[20] ),
    .A2(_04526_),
    .B1(_04537_),
    .B2(\rbzero.spi_registers.texadd2[20] ),
    .X(_04546_));
 sky130_fd_sc_hd__a211o_1 _11355_ (.A1(\rbzero.spi_registers.texadd1[20] ),
    .A2(_04545_),
    .B1(_04536_),
    .C1(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__o21a_1 _11356_ (.A1(\rbzero.spi_registers.texadd0[20] ),
    .A2(_04535_),
    .B1(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__nand2_1 _11357_ (.A(_04544_),
    .B(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__a22o_1 _11358_ (.A1(\rbzero.spi_registers.texadd3[21] ),
    .A2(_04526_),
    .B1(_04537_),
    .B2(\rbzero.spi_registers.texadd2[21] ),
    .X(_04550_));
 sky130_fd_sc_hd__a211o_1 _11359_ (.A1(\rbzero.spi_registers.texadd1[21] ),
    .A2(_04545_),
    .B1(_04536_),
    .C1(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__o21ai_1 _11360_ (.A1(\rbzero.spi_registers.texadd0[21] ),
    .A2(_04535_),
    .B1(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__or3_1 _11361_ (.A(_04454_),
    .B(_04544_),
    .C(_04548_),
    .X(_04553_));
 sky130_fd_sc_hd__a22oi_1 _11362_ (.A1(_04454_),
    .A2(_04552_),
    .B1(_04553_),
    .B2(_04549_),
    .Y(_04554_));
 sky130_fd_sc_hd__a31oi_1 _11363_ (.A1(_04454_),
    .A2(_04549_),
    .A3(_04552_),
    .B1(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__or2_1 _11364_ (.A(\rbzero.spi_registers.texadd0[23] ),
    .B(_04535_),
    .X(_04556_));
 sky130_fd_sc_hd__a22o_1 _11365_ (.A1(\rbzero.spi_registers.texadd3[23] ),
    .A2(_04526_),
    .B1(_04537_),
    .B2(\rbzero.spi_registers.texadd2[23] ),
    .X(_04557_));
 sky130_fd_sc_hd__a211o_1 _11366_ (.A1(\rbzero.spi_registers.texadd1[23] ),
    .A2(_04545_),
    .B1(_04536_),
    .C1(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__a21o_1 _11367_ (.A1(_04556_),
    .A2(_04558_),
    .B1(_03970_),
    .X(_04559_));
 sky130_fd_sc_hd__a221o_1 _11368_ (.A1(\rbzero.spi_registers.texadd2[22] ),
    .A2(\rbzero.wall_hot[0] ),
    .B1(_04545_),
    .B2(\rbzero.spi_registers.texadd1[22] ),
    .C1(_04536_),
    .X(_04560_));
 sky130_fd_sc_hd__a21o_1 _11369_ (.A1(\rbzero.spi_registers.texadd3[22] ),
    .A2(_04526_),
    .B1(_04560_),
    .X(_04561_));
 sky130_fd_sc_hd__o21ai_1 _11370_ (.A1(\rbzero.spi_registers.texadd0[22] ),
    .A2(_04535_),
    .B1(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__nand2_1 _11371_ (.A(_03970_),
    .B(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__or2_1 _11372_ (.A(_04549_),
    .B(_04552_),
    .X(_04564_));
 sky130_fd_sc_hd__mux2_1 _11373_ (.A0(_04562_),
    .A1(_04563_),
    .S(_04564_),
    .X(_04565_));
 sky130_fd_sc_hd__xnor2_1 _11374_ (.A(_04559_),
    .B(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__mux2_1 _11375_ (.A0(_04555_),
    .A1(_04566_),
    .S(_04449_),
    .X(_04567_));
 sky130_fd_sc_hd__or2_1 _11376_ (.A(_04452_),
    .B(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__or3_1 _11377_ (.A(_04454_),
    .B(_04534_),
    .C(_04540_),
    .X(_04569_));
 sky130_fd_sc_hd__a21bo_1 _11378_ (.A1(_04534_),
    .A2(_04540_),
    .B1_N(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__o21ai_1 _11379_ (.A1(_03971_),
    .A2(_04543_),
    .B1(_04570_),
    .Y(_04571_));
 sky130_fd_sc_hd__a211o_1 _11380_ (.A1(_04534_),
    .A2(_04540_),
    .B1(_04543_),
    .C1(_03971_),
    .X(_04572_));
 sky130_fd_sc_hd__and3_1 _11381_ (.A(_03970_),
    .B(_04525_),
    .C(_04529_),
    .X(_04573_));
 sky130_fd_sc_hd__o22ai_1 _11382_ (.A1(_03971_),
    .A2(_04533_),
    .B1(_04573_),
    .B2(_04530_),
    .Y(_04574_));
 sky130_fd_sc_hd__buf_4 _11383_ (.A(\gpout0.hpos[1] ),
    .X(_04575_));
 sky130_fd_sc_hd__o311a_1 _11384_ (.A1(_03971_),
    .A2(_04530_),
    .A3(_04533_),
    .B1(_04574_),
    .C1(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__a311o_1 _11385_ (.A1(_04449_),
    .A2(_04571_),
    .A3(_04572_),
    .B1(_04576_),
    .C1(_04446_),
    .X(_04577_));
 sky130_fd_sc_hd__clkbuf_4 _11386_ (.A(\gpout0.hpos[4] ),
    .X(_04578_));
 sky130_fd_sc_hd__or2_1 _11387_ (.A(_04412_),
    .B(_04578_),
    .X(_04579_));
 sky130_fd_sc_hd__a31o_1 _11388_ (.A1(_04419_),
    .A2(_04568_),
    .A3(_04577_),
    .B1(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__or3_1 _11389_ (.A(_04458_),
    .B(_04521_),
    .C(_04524_),
    .X(_04581_));
 sky130_fd_sc_hd__nor2_1 _11390_ (.A(_04449_),
    .B(_04517_),
    .Y(_04582_));
 sky130_fd_sc_hd__o31a_1 _11391_ (.A1(_04473_),
    .A2(_04513_),
    .A3(_04516_),
    .B1(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__a311oi_2 _11392_ (.A1(_04449_),
    .A2(_04581_),
    .A3(_04525_),
    .B1(_04583_),
    .C1(_03971_),
    .Y(_04584_));
 sky130_fd_sc_hd__a211oi_1 _11393_ (.A1(_04518_),
    .A2(_04520_),
    .B1(_04462_),
    .C1(_04517_),
    .Y(_04585_));
 sky130_fd_sc_hd__and3_1 _11394_ (.A(_04512_),
    .B(_04477_),
    .C(_04510_),
    .X(_04586_));
 sky130_fd_sc_hd__or3_1 _11395_ (.A(_04449_),
    .B(_04513_),
    .C(_04586_),
    .X(_04587_));
 sky130_fd_sc_hd__o311a_1 _11396_ (.A1(_04575_),
    .A2(_04521_),
    .A3(_04585_),
    .B1(_04587_),
    .C1(_03971_),
    .X(_04588_));
 sky130_fd_sc_hd__clkbuf_4 _11397_ (.A(_04578_),
    .X(_04589_));
 sky130_fd_sc_hd__and3_1 _11398_ (.A(_04509_),
    .B(_04481_),
    .C(_04507_),
    .X(_04590_));
 sky130_fd_sc_hd__nand2_1 _11399_ (.A(_04454_),
    .B(_04510_),
    .Y(_04591_));
 sky130_fd_sc_hd__nand2_1 _11400_ (.A(_03970_),
    .B(_04507_),
    .Y(_04592_));
 sky130_fd_sc_hd__a31o_1 _11401_ (.A1(_04506_),
    .A2(_04485_),
    .A3(_04504_),
    .B1(_04592_),
    .X(_04593_));
 sky130_fd_sc_hd__o21ai_1 _11402_ (.A1(_04590_),
    .A2(_04591_),
    .B1(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__nand2_1 _11403_ (.A(_04454_),
    .B(_04504_),
    .Y(_04595_));
 sky130_fd_sc_hd__a21oi_1 _11404_ (.A1(_04501_),
    .A2(_04503_),
    .B1(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__xnor2_1 _11405_ (.A(_04489_),
    .B(_04499_),
    .Y(_04597_));
 sky130_fd_sc_hd__a21o_1 _11406_ (.A1(_03970_),
    .A2(_04597_),
    .B1(_04449_),
    .X(_04598_));
 sky130_fd_sc_hd__o221a_1 _11407_ (.A1(_04575_),
    .A2(_04594_),
    .B1(_04596_),
    .B2(_04598_),
    .C1(_04452_),
    .X(_04599_));
 sky130_fd_sc_hd__nor2_1 _11408_ (.A(_04589_),
    .B(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__o31ai_1 _11409_ (.A1(_04452_),
    .A2(_04584_),
    .A3(_04588_),
    .B1(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__a21o_1 _11410_ (.A1(_04494_),
    .A2(_04495_),
    .B1(\rbzero.texu_hot[0] ),
    .X(_04602_));
 sky130_fd_sc_hd__and2_1 _11411_ (.A(_04496_),
    .B(_04602_),
    .X(_04603_));
 sky130_fd_sc_hd__nand2_1 _11412_ (.A(_04496_),
    .B(_04497_),
    .Y(_04604_));
 sky130_fd_sc_hd__nor2_1 _11413_ (.A(_03970_),
    .B(_04498_),
    .Y(_04605_));
 sky130_fd_sc_hd__a221o_1 _11414_ (.A1(_03970_),
    .A2(_04603_),
    .B1(_04604_),
    .B2(_04605_),
    .C1(_04575_),
    .X(_04606_));
 sky130_fd_sc_hd__a22o_1 _11415_ (.A1(\rbzero.spi_registers.texadd2[5] ),
    .A2(_04537_),
    .B1(_04545_),
    .B2(\rbzero.spi_registers.texadd1[5] ),
    .X(_04607_));
 sky130_fd_sc_hd__a221o_1 _11416_ (.A1(\rbzero.spi_registers.texadd3[5] ),
    .A2(_04457_),
    .B1(_04536_),
    .B2(\rbzero.spi_registers.texadd0[5] ),
    .C1(_03970_),
    .X(_04608_));
 sky130_fd_sc_hd__a22o_1 _11417_ (.A1(\rbzero.spi_registers.texadd2[4] ),
    .A2(_04537_),
    .B1(_04545_),
    .B2(\rbzero.spi_registers.texadd1[4] ),
    .X(_04609_));
 sky130_fd_sc_hd__a221o_1 _11418_ (.A1(\rbzero.spi_registers.texadd3[4] ),
    .A2(_04457_),
    .B1(_04536_),
    .B2(\rbzero.spi_registers.texadd0[4] ),
    .C1(_04454_),
    .X(_04610_));
 sky130_fd_sc_hd__or2_1 _11419_ (.A(_04609_),
    .B(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__o21ai_1 _11420_ (.A1(_04607_),
    .A2(_04608_),
    .B1(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hd__a21oi_1 _11421_ (.A1(_04575_),
    .A2(_04612_),
    .B1(_04452_),
    .Y(_04613_));
 sky130_fd_sc_hd__a22o_1 _11422_ (.A1(\rbzero.spi_registers.texadd2[1] ),
    .A2(_04537_),
    .B1(_04457_),
    .B2(\rbzero.spi_registers.texadd3[1] ),
    .X(_04614_));
 sky130_fd_sc_hd__a21o_1 _11423_ (.A1(\rbzero.spi_registers.texadd1[1] ),
    .A2(_04545_),
    .B1(_04536_),
    .X(_04615_));
 sky130_fd_sc_hd__o221a_1 _11424_ (.A1(\rbzero.spi_registers.texadd0[1] ),
    .A2(_04535_),
    .B1(_04614_),
    .B2(_04615_),
    .C1(_04454_),
    .X(_04616_));
 sky130_fd_sc_hd__a22o_1 _11425_ (.A1(\rbzero.spi_registers.texadd2[0] ),
    .A2(_04537_),
    .B1(_04457_),
    .B2(\rbzero.spi_registers.texadd3[0] ),
    .X(_04617_));
 sky130_fd_sc_hd__a211o_1 _11426_ (.A1(\rbzero.spi_registers.texadd1[0] ),
    .A2(_04545_),
    .B1(_04536_),
    .C1(_04617_),
    .X(_04618_));
 sky130_fd_sc_hd__o211a_1 _11427_ (.A1(\rbzero.spi_registers.texadd0[0] ),
    .A2(_04535_),
    .B1(_04618_),
    .C1(_03970_),
    .X(_04619_));
 sky130_fd_sc_hd__a22o_1 _11428_ (.A1(\rbzero.spi_registers.texadd2[2] ),
    .A2(_04537_),
    .B1(_04457_),
    .B2(\rbzero.spi_registers.texadd3[2] ),
    .X(_04620_));
 sky130_fd_sc_hd__a211o_1 _11429_ (.A1(\rbzero.spi_registers.texadd1[2] ),
    .A2(_04545_),
    .B1(_04536_),
    .C1(_04620_),
    .X(_04621_));
 sky130_fd_sc_hd__o211a_1 _11430_ (.A1(\rbzero.spi_registers.texadd0[2] ),
    .A2(_04535_),
    .B1(_04621_),
    .C1(_03969_),
    .X(_04622_));
 sky130_fd_sc_hd__a22o_1 _11431_ (.A1(\rbzero.spi_registers.texadd3[3] ),
    .A2(_04457_),
    .B1(_04545_),
    .B2(\rbzero.spi_registers.texadd1[3] ),
    .X(_04623_));
 sky130_fd_sc_hd__o21a_1 _11432_ (.A1(\rbzero.spi_registers.texadd2[3] ),
    .A2(_04526_),
    .B1(\rbzero.wall_hot[0] ),
    .X(_04624_));
 sky130_fd_sc_hd__o221a_1 _11433_ (.A1(\rbzero.spi_registers.texadd0[3] ),
    .A2(_04535_),
    .B1(_04623_),
    .B2(_04624_),
    .C1(_04454_),
    .X(_04625_));
 sky130_fd_sc_hd__or3_1 _11434_ (.A(_04575_),
    .B(_04622_),
    .C(_04625_),
    .X(_04626_));
 sky130_fd_sc_hd__o311a_1 _11435_ (.A1(_04449_),
    .A2(_04616_),
    .A3(_04619_),
    .B1(_04626_),
    .C1(_04452_),
    .X(_04627_));
 sky130_fd_sc_hd__buf_4 _11436_ (.A(_04412_),
    .X(_04628_));
 sky130_fd_sc_hd__a211o_1 _11437_ (.A1(_04606_),
    .A2(_04613_),
    .B1(_04627_),
    .C1(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__xnor2_2 _11438_ (.A(_04410_),
    .B(_04423_),
    .Y(_04630_));
 sky130_fd_sc_hd__and3_1 _11439_ (.A(_04601_),
    .B(_04629_),
    .C(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__nor2_1 _11440_ (.A(_04628_),
    .B(_04589_),
    .Y(_04632_));
 sky130_fd_sc_hd__o211a_1 _11441_ (.A1(_04631_),
    .A2(_04632_),
    .B1(_04422_),
    .C1(_04426_),
    .X(_04633_));
 sky130_fd_sc_hd__a32o_2 _11442_ (.A1(_04415_),
    .A2(_04426_),
    .A3(_04451_),
    .B1(_04580_),
    .B2(_04633_),
    .X(net72));
 sky130_fd_sc_hd__buf_1 _11443_ (.A(clknet_leaf_35_i_clk),
    .X(_04634_));
 sky130_fd_sc_hd__inv_2 _20567__3 (.A(clknet_1_1__leaf__03457_),
    .Y(net127));
 sky130_fd_sc_hd__clkinv_2 _11445_ (.A(net2),
    .Y(_04635_));
 sky130_fd_sc_hd__nor2_4 _11446_ (.A(_04445_),
    .B(_04448_),
    .Y(_04636_));
 sky130_fd_sc_hd__and2_1 _11447_ (.A(\gpout0.hpos[3] ),
    .B(_04636_),
    .X(_04637_));
 sky130_fd_sc_hd__or2_2 _11448_ (.A(\gpout0.hpos[4] ),
    .B(_04637_),
    .X(_04638_));
 sky130_fd_sc_hd__o21a_1 _11449_ (.A1(\gpout0.hpos[5] ),
    .A2(_04638_),
    .B1(\gpout0.hpos[6] ),
    .X(_04639_));
 sky130_fd_sc_hd__and2_1 _11450_ (.A(\gpout0.hpos[7] ),
    .B(_04639_),
    .X(_04640_));
 sky130_fd_sc_hd__a21oi_2 _11451_ (.A1(\gpout0.hpos[8] ),
    .A2(_04640_),
    .B1(\gpout0.hpos[9] ),
    .Y(_04641_));
 sky130_fd_sc_hd__buf_2 _11452_ (.A(\gpout0.vpos[7] ),
    .X(_04642_));
 sky130_fd_sc_hd__clkinv_4 _11453_ (.A(net3),
    .Y(_04643_));
 sky130_fd_sc_hd__or4_1 _11454_ (.A(\gpout0.vpos[9] ),
    .B(\gpout0.vpos[8] ),
    .C(_04642_),
    .D(_04643_),
    .X(_04644_));
 sky130_fd_sc_hd__or2_1 _11455_ (.A(\gpout0.vpos[5] ),
    .B(\gpout0.vpos[4] ),
    .X(_04645_));
 sky130_fd_sc_hd__or2_1 _11456_ (.A(\gpout0.vpos[3] ),
    .B(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__or3_2 _11457_ (.A(\gpout0.vpos[2] ),
    .B(\gpout0.vpos[1] ),
    .C(\gpout0.vpos[0] ),
    .X(_04647_));
 sky130_fd_sc_hd__clkbuf_4 _11458_ (.A(\gpout0.vpos[6] ),
    .X(_04648_));
 sky130_fd_sc_hd__o21a_1 _11459_ (.A1(_04646_),
    .A2(_04647_),
    .B1(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__nor3_4 _11460_ (.A(_04641_),
    .B(_04644_),
    .C(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__clkbuf_4 _11461_ (.A(\gpout0.vpos[4] ),
    .X(_04651_));
 sky130_fd_sc_hd__buf_4 _11462_ (.A(\gpout0.vpos[3] ),
    .X(_04652_));
 sky130_fd_sc_hd__clkbuf_4 _11463_ (.A(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__or2_1 _11464_ (.A(_04651_),
    .B(_04653_),
    .X(_04654_));
 sky130_fd_sc_hd__nand2_1 _11465_ (.A(_04651_),
    .B(_04652_),
    .Y(_04655_));
 sky130_fd_sc_hd__clkbuf_4 _11466_ (.A(\gpout0.vpos[5] ),
    .X(_04656_));
 sky130_fd_sc_hd__clkbuf_4 _11467_ (.A(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__nand2_1 _11468_ (.A(_04657_),
    .B(_04651_),
    .Y(_04658_));
 sky130_fd_sc_hd__o21ai_1 _11469_ (.A1(_04446_),
    .A2(_04448_),
    .B1(_04647_),
    .Y(_04659_));
 sky130_fd_sc_hd__a41o_1 _11470_ (.A1(_04645_),
    .A2(_04654_),
    .A3(_04655_),
    .A4(_04658_),
    .B1(_04659_),
    .X(_04660_));
 sky130_fd_sc_hd__and2_1 _11471_ (.A(_04650_),
    .B(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__nand2_1 _11472_ (.A(_04656_),
    .B(\rbzero.debug_overlay.playerY[2] ),
    .Y(_04662_));
 sky130_fd_sc_hd__or2_1 _11473_ (.A(_04656_),
    .B(\rbzero.debug_overlay.playerY[2] ),
    .X(_04663_));
 sky130_fd_sc_hd__nand2_1 _11474_ (.A(_04653_),
    .B(\rbzero.debug_overlay.playerY[0] ),
    .Y(_04664_));
 sky130_fd_sc_hd__or2_1 _11475_ (.A(_04652_),
    .B(\rbzero.debug_overlay.playerY[0] ),
    .X(_04665_));
 sky130_fd_sc_hd__a22o_1 _11476_ (.A1(_04662_),
    .A2(_04663_),
    .B1(_04664_),
    .B2(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__inv_2 _11477_ (.A(\rbzero.debug_overlay.playerY[3] ),
    .Y(_04667_));
 sky130_fd_sc_hd__xnor2_1 _11478_ (.A(_04651_),
    .B(\rbzero.debug_overlay.playerY[1] ),
    .Y(_04668_));
 sky130_fd_sc_hd__o221a_1 _11479_ (.A1(_04648_),
    .A2(_04667_),
    .B1(\rbzero.debug_overlay.playerX[0] ),
    .B2(_04413_),
    .C1(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__clkinv_2 _11480_ (.A(\gpout0.vpos[7] ),
    .Y(_04670_));
 sky130_fd_sc_hd__inv_2 _11481_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .Y(_04671_));
 sky130_fd_sc_hd__inv_2 _11482_ (.A(\gpout0.vpos[6] ),
    .Y(_04672_));
 sky130_fd_sc_hd__inv_2 _11483_ (.A(\rbzero.debug_overlay.playerY[4] ),
    .Y(_04673_));
 sky130_fd_sc_hd__clkinv_2 _11484_ (.A(\rbzero.debug_overlay.playerX[2] ),
    .Y(_04674_));
 sky130_fd_sc_hd__o22a_1 _11485_ (.A1(\gpout0.vpos[7] ),
    .A2(_04673_),
    .B1(_04674_),
    .B2(_04411_),
    .X(_04675_));
 sky130_fd_sc_hd__o221a_1 _11486_ (.A1(_04672_),
    .A2(\rbzero.debug_overlay.playerY[3] ),
    .B1(\rbzero.debug_overlay.playerX[2] ),
    .B2(_04421_),
    .C1(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__o221a_1 _11487_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_04410_),
    .B1(_04578_),
    .B2(_04671_),
    .C1(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__o221a_1 _11488_ (.A1(_04670_),
    .A2(\rbzero.debug_overlay.playerY[4] ),
    .B1(\rbzero.debug_overlay.playerX[1] ),
    .B2(_04414_),
    .C1(_04677_),
    .X(_04678_));
 sky130_fd_sc_hd__inv_2 _11489_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .Y(_04679_));
 sky130_fd_sc_hd__inv_2 _11490_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .Y(_04680_));
 sky130_fd_sc_hd__xnor2_1 _11491_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .B(_03972_),
    .Y(_04681_));
 sky130_fd_sc_hd__o221a_1 _11492_ (.A1(_04679_),
    .A2(_04628_),
    .B1(_04419_),
    .B2(_04680_),
    .C1(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__and4b_1 _11493_ (.A_N(_04666_),
    .B(_04669_),
    .C(_04678_),
    .D(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__xnor2_1 _11494_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_03969_),
    .Y(_04684_));
 sky130_fd_sc_hd__xnor2_1 _11495_ (.A(\gpout0.vpos[1] ),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .Y(_04685_));
 sky130_fd_sc_hd__inv_2 _11496_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .Y(_04686_));
 sky130_fd_sc_hd__clkbuf_4 _11497_ (.A(\gpout0.vpos[2] ),
    .X(_04687_));
 sky130_fd_sc_hd__xnor2_1 _11498_ (.A(_04687_),
    .B(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_04688_));
 sky130_fd_sc_hd__o221a_1 _11499_ (.A1(\gpout0.vpos[0] ),
    .A2(_04686_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .B2(_04446_),
    .C1(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__and3_1 _11500_ (.A(_04684_),
    .B(_04685_),
    .C(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__inv_2 _11501_ (.A(\gpout0.vpos[0] ),
    .Y(_04691_));
 sky130_fd_sc_hd__inv_2 _11502_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .Y(_04692_));
 sky130_fd_sc_hd__xnor2_1 _11503_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(\gpout0.hpos[1] ),
    .Y(_04693_));
 sky130_fd_sc_hd__o221a_1 _11504_ (.A1(_04691_),
    .A2(\rbzero.debug_overlay.playerY[-3] ),
    .B1(_04692_),
    .B2(\gpout0.hpos[2] ),
    .C1(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__or3_1 _11505_ (.A(_04642_),
    .B(_04648_),
    .C(_04645_),
    .X(_04695_));
 sky130_fd_sc_hd__o31a_1 _11506_ (.A1(_04653_),
    .A2(_04647_),
    .A3(_04695_),
    .B1(\gpout0.vpos[8] ),
    .X(_04696_));
 sky130_fd_sc_hd__or3b_1 _11507_ (.A(\gpout0.vpos[9] ),
    .B(_04420_),
    .C_N(net1),
    .X(_04697_));
 sky130_fd_sc_hd__or2_1 _11508_ (.A(\gpout0.hpos[2] ),
    .B(_04447_),
    .X(_04698_));
 sky130_fd_sc_hd__or2_1 _11509_ (.A(\gpout0.hpos[6] ),
    .B(\gpout0.hpos[5] ),
    .X(_04699_));
 sky130_fd_sc_hd__or2_1 _11510_ (.A(_04579_),
    .B(_04699_),
    .X(_04700_));
 sky130_fd_sc_hd__o31a_1 _11511_ (.A1(_03972_),
    .A2(_04698_),
    .A3(_04700_),
    .B1(\gpout0.hpos[8] ),
    .X(_04701_));
 sky130_fd_sc_hd__or3_2 _11512_ (.A(_04696_),
    .B(_04697_),
    .C(_04701_),
    .X(_04702_));
 sky130_fd_sc_hd__a31o_1 _11513_ (.A1(_04683_),
    .A2(_04690_),
    .A3(_04694_),
    .B1(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__buf_4 _11514_ (.A(_04411_),
    .X(_04704_));
 sky130_fd_sc_hd__inv_2 _11515_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .Y(_04705_));
 sky130_fd_sc_hd__xor2_1 _11516_ (.A(\gpout0.vpos[4] ),
    .B(\rbzero.map_overlay.i_othery[1] ),
    .X(_04706_));
 sky130_fd_sc_hd__a221o_1 _11517_ (.A1(\rbzero.map_overlay.i_otherx[3] ),
    .A2(_04410_),
    .B1(_04704_),
    .B2(_04705_),
    .C1(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__inv_2 _11518_ (.A(\rbzero.map_overlay.i_otherx[1] ),
    .Y(_04708_));
 sky130_fd_sc_hd__xnor2_1 _11519_ (.A(_04656_),
    .B(\rbzero.map_overlay.i_othery[2] ),
    .Y(_04709_));
 sky130_fd_sc_hd__o221a_1 _11520_ (.A1(_04670_),
    .A2(\rbzero.map_overlay.i_othery[4] ),
    .B1(_04708_),
    .B2(_04578_),
    .C1(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__xnor2_1 _11521_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .B(_03972_),
    .Y(_04711_));
 sky130_fd_sc_hd__xnor2_1 _11522_ (.A(_04652_),
    .B(\rbzero.map_overlay.i_othery[0] ),
    .Y(_04712_));
 sky130_fd_sc_hd__inv_2 _11523_ (.A(\rbzero.map_overlay.i_othery[4] ),
    .Y(_04713_));
 sky130_fd_sc_hd__xnor2_1 _11524_ (.A(_04648_),
    .B(\rbzero.map_overlay.i_othery[3] ),
    .Y(_04714_));
 sky130_fd_sc_hd__o221a_1 _11525_ (.A1(\gpout0.vpos[7] ),
    .A2(_04713_),
    .B1(\rbzero.map_overlay.i_otherx[1] ),
    .B2(_04414_),
    .C1(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__xnor2_1 _11526_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .B(_04412_),
    .Y(_04716_));
 sky130_fd_sc_hd__o221a_1 _11527_ (.A1(\rbzero.map_overlay.i_otherx[3] ),
    .A2(_04410_),
    .B1(_04411_),
    .B2(_04705_),
    .C1(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__and4_1 _11528_ (.A(_04711_),
    .B(_04712_),
    .C(_04715_),
    .D(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__and3b_1 _11529_ (.A_N(_04707_),
    .B(_04710_),
    .C(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__inv_2 _11530_ (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .Y(_04720_));
 sky130_fd_sc_hd__inv_2 _11531_ (.A(\rbzero.map_overlay.i_mapdx[1] ),
    .Y(_04721_));
 sky130_fd_sc_hd__a22o_1 _11532_ (.A1(_04720_),
    .A2(_03973_),
    .B1(_04578_),
    .B2(_04721_),
    .X(_04722_));
 sky130_fd_sc_hd__xor2_1 _11533_ (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(_04704_),
    .X(_04723_));
 sky130_fd_sc_hd__a22o_1 _11534_ (.A1(\rbzero.map_overlay.i_mapdx[0] ),
    .A2(_04413_),
    .B1(_04414_),
    .B2(\rbzero.map_overlay.i_mapdx[1] ),
    .X(_04724_));
 sky130_fd_sc_hd__or4_1 _11535_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(\rbzero.map_overlay.i_mapdx[2] ),
    .C(\rbzero.map_overlay.i_mapdx[1] ),
    .D(\rbzero.map_overlay.i_mapdx[0] ),
    .X(_04725_));
 sky130_fd_sc_hd__o21a_1 _11536_ (.A1(\rbzero.map_overlay.i_mapdx[5] ),
    .A2(_04725_),
    .B1(_04720_),
    .X(_04726_));
 sky130_fd_sc_hd__xnor2_1 _11537_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_04418_),
    .Y(_04727_));
 sky130_fd_sc_hd__o221a_1 _11538_ (.A1(\rbzero.map_overlay.i_mapdx[0] ),
    .A2(_04413_),
    .B1(_03972_),
    .B2(_04726_),
    .C1(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__or3b_1 _11539_ (.A(_04723_),
    .B(_04724_),
    .C_N(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__inv_2 _11540_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .Y(_04730_));
 sky130_fd_sc_hd__inv_2 _11541_ (.A(_04656_),
    .Y(_04731_));
 sky130_fd_sc_hd__xnor2_1 _11542_ (.A(_04651_),
    .B(\rbzero.map_overlay.i_mapdy[1] ),
    .Y(_04732_));
 sky130_fd_sc_hd__o221a_1 _11543_ (.A1(_04648_),
    .A2(_04730_),
    .B1(\rbzero.map_overlay.i_mapdy[2] ),
    .B2(_04731_),
    .C1(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__a22oi_1 _11544_ (.A1(_04670_),
    .A2(\rbzero.map_overlay.i_mapdy[4] ),
    .B1(\rbzero.map_overlay.i_mapdy[2] ),
    .B2(_04731_),
    .Y(_04734_));
 sky130_fd_sc_hd__inv_2 _11545_ (.A(_04652_),
    .Y(_04735_));
 sky130_fd_sc_hd__or4_1 _11546_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(\rbzero.map_overlay.i_mapdy[2] ),
    .C(\rbzero.map_overlay.i_mapdy[1] ),
    .D(\rbzero.map_overlay.i_mapdy[0] ),
    .X(_04736_));
 sky130_fd_sc_hd__o21a_1 _11547_ (.A1(\rbzero.map_overlay.i_mapdy[5] ),
    .A2(_04736_),
    .B1(_04670_),
    .X(_04737_));
 sky130_fd_sc_hd__inv_2 _11548_ (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .Y(_04738_));
 sky130_fd_sc_hd__o22a_1 _11549_ (.A1(_04672_),
    .A2(\rbzero.map_overlay.i_mapdy[3] ),
    .B1(_04738_),
    .B2(_04653_),
    .X(_04739_));
 sky130_fd_sc_hd__o221a_1 _11550_ (.A1(_04735_),
    .A2(\rbzero.map_overlay.i_mapdy[0] ),
    .B1(_04737_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_04739_),
    .X(_04740_));
 sky130_fd_sc_hd__and3_1 _11551_ (.A(_04733_),
    .B(_04734_),
    .C(_04740_),
    .X(_04741_));
 sky130_fd_sc_hd__o21a_1 _11552_ (.A1(_04722_),
    .A2(_04729_),
    .B1(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__nand2_1 _11553_ (.A(_04698_),
    .B(_04647_),
    .Y(_04743_));
 sky130_fd_sc_hd__nor2_1 _11554_ (.A(_04683_),
    .B(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__o21a_1 _11555_ (.A1(_04719_),
    .A2(_04742_),
    .B1(_04744_),
    .X(_04745_));
 sky130_fd_sc_hd__nand2_1 _11556_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_04746_));
 sky130_fd_sc_hd__or2_1 _11557_ (.A(\rbzero.traced_texVinit[9] ),
    .B(\rbzero.texV[9] ),
    .X(_04747_));
 sky130_fd_sc_hd__and2_1 _11558_ (.A(_04746_),
    .B(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__nand2_1 _11559_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .Y(_04749_));
 sky130_fd_sc_hd__or2_1 _11560_ (.A(\rbzero.traced_texVinit[8] ),
    .B(\rbzero.spi_registers.vshift[5] ),
    .X(_04750_));
 sky130_fd_sc_hd__and3_1 _11561_ (.A(\rbzero.texV[8] ),
    .B(_04749_),
    .C(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__a21o_1 _11562_ (.A1(\rbzero.traced_texVinit[8] ),
    .A2(\rbzero.spi_registers.vshift[5] ),
    .B1(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__nand2_1 _11563_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .Y(_04753_));
 sky130_fd_sc_hd__or2_1 _11564_ (.A(\rbzero.traced_texVinit[7] ),
    .B(\rbzero.spi_registers.vshift[4] ),
    .X(_04754_));
 sky130_fd_sc_hd__nand2_1 _11565_ (.A(_04753_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__xor2_1 _11566_ (.A(\rbzero.texV[7] ),
    .B(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__nand2_1 _11567_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .Y(_04757_));
 sky130_fd_sc_hd__or2_1 _11568_ (.A(\rbzero.traced_texVinit[6] ),
    .B(\rbzero.spi_registers.vshift[3] ),
    .X(_04758_));
 sky130_fd_sc_hd__nand3_1 _11569_ (.A(\rbzero.texV[6] ),
    .B(_04757_),
    .C(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__nand3_1 _11570_ (.A(_04756_),
    .B(_04757_),
    .C(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__a21o_1 _11571_ (.A1(_04757_),
    .A2(_04758_),
    .B1(\rbzero.texV[6] ),
    .X(_04761_));
 sky130_fd_sc_hd__nand2_1 _11572_ (.A(_04759_),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__and2_1 _11573_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .X(_04763_));
 sky130_fd_sc_hd__nor2_1 _11574_ (.A(\rbzero.traced_texVinit[5] ),
    .B(\rbzero.spi_registers.vshift[2] ),
    .Y(_04764_));
 sky130_fd_sc_hd__nor2_1 _11575_ (.A(_04763_),
    .B(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__a21oi_2 _11576_ (.A1(\rbzero.texV[5] ),
    .A2(_04765_),
    .B1(_04763_),
    .Y(_04766_));
 sky130_fd_sc_hd__xnor2_1 _11577_ (.A(_04762_),
    .B(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__nand2_1 _11578_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .Y(_04768_));
 sky130_fd_sc_hd__or2_1 _11579_ (.A(\rbzero.traced_texVinit[4] ),
    .B(\rbzero.spi_registers.vshift[1] ),
    .X(_04769_));
 sky130_fd_sc_hd__nand3_1 _11580_ (.A(\rbzero.texV[4] ),
    .B(_04768_),
    .C(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hd__xnor2_1 _11581_ (.A(\rbzero.texV[5] ),
    .B(_04765_),
    .Y(_04771_));
 sky130_fd_sc_hd__a21oi_1 _11582_ (.A1(_04768_),
    .A2(_04770_),
    .B1(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__a21o_1 _11583_ (.A1(_04768_),
    .A2(_04769_),
    .B1(\rbzero.texV[4] ),
    .X(_04773_));
 sky130_fd_sc_hd__nand2_1 _11584_ (.A(_04770_),
    .B(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__or2_1 _11585_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .X(_04775_));
 sky130_fd_sc_hd__nand2_1 _11586_ (.A(\rbzero.traced_texVinit[3] ),
    .B(\rbzero.spi_registers.vshift[0] ),
    .Y(_04776_));
 sky130_fd_sc_hd__a21boi_1 _11587_ (.A1(\rbzero.texV[3] ),
    .A2(_04775_),
    .B1_N(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__nor2_1 _11588_ (.A(_04774_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__xnor2_1 _11589_ (.A(_04774_),
    .B(_04777_),
    .Y(_04779_));
 sky130_fd_sc_hd__nand2_1 _11590_ (.A(_04776_),
    .B(_04775_),
    .Y(_04780_));
 sky130_fd_sc_hd__xor2_2 _11591_ (.A(\rbzero.texV[3] ),
    .B(_04780_),
    .X(_04781_));
 sky130_fd_sc_hd__o211a_1 _11592_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(\rbzero.texV[1] ),
    .B1(\rbzero.texV[0] ),
    .C1(\rbzero.traced_texVinit[0] ),
    .X(_04782_));
 sky130_fd_sc_hd__a221o_1 _11593_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(\rbzero.texV[1] ),
    .B2(\rbzero.traced_texVinit[1] ),
    .C1(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__o21ai_2 _11594_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(\rbzero.texV[2] ),
    .B1(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__or2_4 _11595_ (.A(_04781_),
    .B(_04784_),
    .X(_04785_));
 sky130_fd_sc_hd__nor2_2 _11596_ (.A(_04779_),
    .B(_04785_),
    .Y(_04786_));
 sky130_fd_sc_hd__and3_1 _11597_ (.A(_04771_),
    .B(_04768_),
    .C(_04770_),
    .X(_04787_));
 sky130_fd_sc_hd__or2_1 _11598_ (.A(_04772_),
    .B(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__inv_2 _11599_ (.A(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__o21a_1 _11600_ (.A1(_04778_),
    .A2(_04786_),
    .B1(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__nor2_1 _11601_ (.A(_04772_),
    .B(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__nor2_1 _11602_ (.A(_04767_),
    .B(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__o21bai_4 _11603_ (.A1(_04762_),
    .A2(_04766_),
    .B1_N(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__a21oi_1 _11604_ (.A1(_04757_),
    .A2(_04759_),
    .B1(_04756_),
    .Y(_04794_));
 sky130_fd_sc_hd__a21o_1 _11605_ (.A1(_04760_),
    .A2(_04793_),
    .B1(_04794_),
    .X(_04795_));
 sky130_fd_sc_hd__a21oi_1 _11606_ (.A1(_04749_),
    .A2(_04750_),
    .B1(\rbzero.texV[8] ),
    .Y(_04796_));
 sky130_fd_sc_hd__a21boi_1 _11607_ (.A1(\rbzero.texV[7] ),
    .A2(_04754_),
    .B1_N(_04753_),
    .Y(_04797_));
 sky130_fd_sc_hd__or3_1 _11608_ (.A(_04751_),
    .B(_04796_),
    .C(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__inv_2 _11609_ (.A(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__o21ai_1 _11610_ (.A1(_04751_),
    .A2(_04796_),
    .B1(_04797_),
    .Y(_04800_));
 sky130_fd_sc_hd__o221a_1 _11611_ (.A1(_04748_),
    .A2(_04752_),
    .B1(_04795_),
    .B2(_04799_),
    .C1(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__a21o_1 _11612_ (.A1(_04748_),
    .A2(_04752_),
    .B1(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__xor2_1 _11613_ (.A(\rbzero.traced_texVinit[10] ),
    .B(\rbzero.texV[10] ),
    .X(_04803_));
 sky130_fd_sc_hd__xnor2_1 _11614_ (.A(_04746_),
    .B(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__a21oi_1 _11615_ (.A1(_04802_),
    .A2(_04804_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_04805_));
 sky130_fd_sc_hd__o21a_4 _11616_ (.A1(_04802_),
    .A2(_04804_),
    .B1(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__and3_1 _11617_ (.A(_04795_),
    .B(_04798_),
    .C(_04800_),
    .X(_04807_));
 sky130_fd_sc_hd__a21o_1 _11618_ (.A1(_04798_),
    .A2(_04800_),
    .B1(_04795_),
    .X(_04808_));
 sky130_fd_sc_hd__or3b_1 _11619_ (.A(_04806_),
    .B(_04807_),
    .C_N(_04808_),
    .X(_04809_));
 sky130_fd_sc_hd__buf_8 _11620_ (.A(_04809_),
    .X(_04810_));
 sky130_fd_sc_hd__and2_1 _11621_ (.A(_04767_),
    .B(_04791_),
    .X(_04811_));
 sky130_fd_sc_hd__nor3_4 _11622_ (.A(_04792_),
    .B(_04806_),
    .C(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__nor3_2 _11623_ (.A(_04789_),
    .B(_04778_),
    .C(_04786_),
    .Y(_04813_));
 sky130_fd_sc_hd__or3_4 _11624_ (.A(_04790_),
    .B(_04806_),
    .C(_04813_),
    .X(_04814_));
 sky130_fd_sc_hd__nand2_1 _11625_ (.A(_04779_),
    .B(_04785_),
    .Y(_04815_));
 sky130_fd_sc_hd__or3b_1 _11626_ (.A(_04786_),
    .B(_04806_),
    .C_N(_04815_),
    .X(_04816_));
 sky130_fd_sc_hd__buf_4 _11627_ (.A(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__nand2_1 _11628_ (.A(_04814_),
    .B(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__or2_1 _11629_ (.A(_04812_),
    .B(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__inv_2 _11630_ (.A(_04760_),
    .Y(_04820_));
 sky130_fd_sc_hd__nor2_2 _11631_ (.A(_04820_),
    .B(_04794_),
    .Y(_04821_));
 sky130_fd_sc_hd__xnor2_4 _11632_ (.A(_04793_),
    .B(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__nor2_8 _11633_ (.A(_04806_),
    .B(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__or2_1 _11634_ (.A(_03972_),
    .B(_04418_),
    .X(_04824_));
 sky130_fd_sc_hd__a21oi_4 _11635_ (.A1(\gpout0.hpos[8] ),
    .A2(_04824_),
    .B1(_04420_),
    .Y(_04825_));
 sky130_fd_sc_hd__nor3b_4 _11636_ (.A(_04786_),
    .B(_04806_),
    .C_N(_04815_),
    .Y(_04826_));
 sky130_fd_sc_hd__buf_4 _11637_ (.A(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__a21oi_4 _11638_ (.A1(_04781_),
    .A2(_04784_),
    .B1(_04806_),
    .Y(_04828_));
 sky130_fd_sc_hd__and2_2 _11639_ (.A(_04785_),
    .B(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__buf_2 _11640_ (.A(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__clkbuf_4 _11641_ (.A(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__inv_4 _11642_ (.A(_04810_),
    .Y(_04832_));
 sky130_fd_sc_hd__or3_1 _11643_ (.A(_04827_),
    .B(_04831_),
    .C(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__or4_1 _11644_ (.A(_04819_),
    .B(_04823_),
    .C(_04825_),
    .D(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__inv_2 _11645_ (.A(\rbzero.row_render.size[2] ),
    .Y(_04835_));
 sky130_fd_sc_hd__nor2_1 _11646_ (.A(\rbzero.row_render.size[1] ),
    .B(\rbzero.row_render.size[0] ),
    .Y(_04836_));
 sky130_fd_sc_hd__nand2_1 _11647_ (.A(_04835_),
    .B(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hd__or2_1 _11648_ (.A(\rbzero.row_render.size[3] ),
    .B(_04837_),
    .X(_04838_));
 sky130_fd_sc_hd__or3_1 _11649_ (.A(\rbzero.row_render.size[5] ),
    .B(\rbzero.row_render.size[4] ),
    .C(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__and2_1 _11650_ (.A(\rbzero.row_render.size[6] ),
    .B(_04839_),
    .X(_04840_));
 sky130_fd_sc_hd__o21a_1 _11651_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_04840_),
    .B1(\rbzero.row_render.size[8] ),
    .X(_04841_));
 sky130_fd_sc_hd__nor3_1 _11652_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(_04840_),
    .Y(_04842_));
 sky130_fd_sc_hd__nor2_1 _11653_ (.A(_04841_),
    .B(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__xnor2_1 _11654_ (.A(\rbzero.row_render.size[7] ),
    .B(_04840_),
    .Y(_04844_));
 sky130_fd_sc_hd__a22o_1 _11655_ (.A1(\gpout0.hpos[7] ),
    .A2(_04844_),
    .B1(_04843_),
    .B2(\gpout0.hpos[8] ),
    .X(_04845_));
 sky130_fd_sc_hd__nor2_1 _11656_ (.A(\rbzero.row_render.size[6] ),
    .B(_04839_),
    .Y(_04846_));
 sky130_fd_sc_hd__nor2_1 _11657_ (.A(_04840_),
    .B(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__o21ai_1 _11658_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_04838_),
    .B1(\rbzero.row_render.size[5] ),
    .Y(_04848_));
 sky130_fd_sc_hd__nand2_1 _11659_ (.A(_04839_),
    .B(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__xnor2_1 _11660_ (.A(\rbzero.row_render.size[4] ),
    .B(_04838_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand2_1 _11661_ (.A(\rbzero.row_render.size[3] ),
    .B(_04837_),
    .Y(_04851_));
 sky130_fd_sc_hd__nand2_1 _11662_ (.A(_04838_),
    .B(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__or2_1 _11663_ (.A(_04835_),
    .B(_04836_),
    .X(_04853_));
 sky130_fd_sc_hd__nor2_1 _11664_ (.A(_04412_),
    .B(_04852_),
    .Y(_04854_));
 sky130_fd_sc_hd__o211a_1 _11665_ (.A1(\rbzero.row_render.size[0] ),
    .A2(\gpout0.hpos[1] ),
    .B1(_04447_),
    .C1(\rbzero.row_render.size[1] ),
    .X(_04855_));
 sky130_fd_sc_hd__a211o_1 _11666_ (.A1(\gpout0.hpos[1] ),
    .A2(_03969_),
    .B1(_04836_),
    .C1(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__a21oi_1 _11667_ (.A1(\rbzero.row_render.size[2] ),
    .A2(\gpout0.hpos[2] ),
    .B1(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__a311oi_1 _11668_ (.A1(_04446_),
    .A2(_04837_),
    .A3(_04853_),
    .B1(_04854_),
    .C1(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__a221o_1 _11669_ (.A1(_04412_),
    .A2(_04852_),
    .B1(_04850_),
    .B2(\gpout0.hpos[4] ),
    .C1(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__o221a_1 _11670_ (.A1(\gpout0.hpos[4] ),
    .A2(_04850_),
    .B1(_04849_),
    .B2(_04411_),
    .C1(_04859_),
    .X(_04860_));
 sky130_fd_sc_hd__a221o_1 _11671_ (.A1(_04411_),
    .A2(_04849_),
    .B1(_04847_),
    .B2(_04418_),
    .C1(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__o221a_1 _11672_ (.A1(_04418_),
    .A2(_04847_),
    .B1(_04844_),
    .B2(\gpout0.hpos[7] ),
    .C1(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__o22a_1 _11673_ (.A1(\gpout0.hpos[8] ),
    .A2(_04843_),
    .B1(_04845_),
    .B2(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__a21o_1 _11674_ (.A1(\rbzero.row_render.size[7] ),
    .A2(\rbzero.row_render.size[6] ),
    .B1(\rbzero.row_render.size[8] ),
    .X(_04864_));
 sky130_fd_sc_hd__nand3_1 _11675_ (.A(\rbzero.row_render.size[8] ),
    .B(\rbzero.row_render.size[7] ),
    .C(\rbzero.row_render.size[6] ),
    .Y(_04865_));
 sky130_fd_sc_hd__a21o_1 _11676_ (.A1(_04864_),
    .A2(_04865_),
    .B1(\gpout0.hpos[8] ),
    .X(_04866_));
 sky130_fd_sc_hd__xnor2_1 _11677_ (.A(\rbzero.row_render.size[7] ),
    .B(\rbzero.row_render.size[6] ),
    .Y(_04867_));
 sky130_fd_sc_hd__o22a_1 _11678_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_04418_),
    .B1(_04867_),
    .B2(\gpout0.hpos[7] ),
    .X(_04868_));
 sky130_fd_sc_hd__and2_1 _11679_ (.A(\rbzero.row_render.size[1] ),
    .B(_04449_),
    .X(_04869_));
 sky130_fd_sc_hd__o22a_1 _11680_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_04446_),
    .B1(_04449_),
    .B2(\rbzero.row_render.size[1] ),
    .X(_04870_));
 sky130_fd_sc_hd__o31a_1 _11681_ (.A1(\rbzero.row_render.size[0] ),
    .A2(_04453_),
    .A3(_04869_),
    .B1(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__a221o_1 _11682_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_04413_),
    .B1(_04446_),
    .B2(\rbzero.row_render.size[2] ),
    .C1(_04871_),
    .X(_04872_));
 sky130_fd_sc_hd__o221a_1 _11683_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_04413_),
    .B1(_04414_),
    .B2(\rbzero.row_render.size[4] ),
    .C1(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__a221o_1 _11684_ (.A1(\rbzero.row_render.size[5] ),
    .A2(_04421_),
    .B1(_04414_),
    .B2(\rbzero.row_render.size[4] ),
    .C1(_04873_),
    .X(_04874_));
 sky130_fd_sc_hd__o2bb2a_1 _11685_ (.A1_N(\rbzero.row_render.size[6] ),
    .A2_N(_04418_),
    .B1(_04421_),
    .B2(\rbzero.row_render.size[5] ),
    .X(_04875_));
 sky130_fd_sc_hd__nand2_1 _11686_ (.A(_04874_),
    .B(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__a22o_1 _11687_ (.A1(_03972_),
    .A2(_04867_),
    .B1(_04868_),
    .B2(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__and3_1 _11688_ (.A(\gpout0.hpos[8] ),
    .B(_04864_),
    .C(_04865_),
    .X(_04878_));
 sky130_fd_sc_hd__a21oi_1 _11689_ (.A1(_04866_),
    .A2(_04877_),
    .B1(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hd__a21o_1 _11690_ (.A1(\rbzero.row_render.size[9] ),
    .A2(_04864_),
    .B1(_03976_),
    .X(_04880_));
 sky130_fd_sc_hd__o21a_1 _11691_ (.A1(\rbzero.row_render.size[9] ),
    .A2(_04864_),
    .B1(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__or2_1 _11692_ (.A(_03976_),
    .B(_04864_),
    .X(_04882_));
 sky130_fd_sc_hd__o221a_1 _11693_ (.A1(\gpout0.hpos[9] ),
    .A2(_04863_),
    .B1(_04879_),
    .B2(_04881_),
    .C1(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__or4_2 _11694_ (.A(\rbzero.row_render.size[10] ),
    .B(\rbzero.row_render.size[9] ),
    .C(_04841_),
    .D(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__a21oi_1 _11695_ (.A1(_04834_),
    .A2(_04884_),
    .B1(\rbzero.row_render.vinf ),
    .Y(_04885_));
 sky130_fd_sc_hd__or2_4 _11696_ (.A(_04806_),
    .B(_04822_),
    .X(_04886_));
 sky130_fd_sc_hd__buf_6 _11697_ (.A(_04886_),
    .X(_04887_));
 sky130_fd_sc_hd__or3_1 _11698_ (.A(_04792_),
    .B(_04806_),
    .C(_04811_),
    .X(_04888_));
 sky130_fd_sc_hd__buf_6 _11699_ (.A(_04888_),
    .X(_04889_));
 sky130_fd_sc_hd__buf_4 _11700_ (.A(_04814_),
    .X(_04890_));
 sky130_fd_sc_hd__buf_4 _11701_ (.A(_04817_),
    .X(_04891_));
 sky130_fd_sc_hd__nand2_4 _11702_ (.A(_04785_),
    .B(_04828_),
    .Y(_04892_));
 sky130_fd_sc_hd__buf_6 _11703_ (.A(_04892_),
    .X(_04893_));
 sky130_fd_sc_hd__o211a_1 _11704_ (.A1(\rbzero.floor_leak[1] ),
    .A2(_04817_),
    .B1(_04893_),
    .C1(\rbzero.floor_leak[0] ),
    .X(_04894_));
 sky130_fd_sc_hd__a221o_1 _11705_ (.A1(\rbzero.floor_leak[2] ),
    .A2(_04814_),
    .B1(_04891_),
    .B2(\rbzero.floor_leak[1] ),
    .C1(_04894_),
    .X(_04895_));
 sky130_fd_sc_hd__o221a_1 _11706_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_04889_),
    .B1(_04890_),
    .B2(\rbzero.floor_leak[2] ),
    .C1(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__a221o_1 _11707_ (.A1(\rbzero.floor_leak[3] ),
    .A2(_04889_),
    .B1(_04886_),
    .B2(\rbzero.floor_leak[4] ),
    .C1(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__o221a_1 _11708_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_04810_),
    .B1(_04887_),
    .B2(\rbzero.floor_leak[4] ),
    .C1(_04897_),
    .X(_04898_));
 sky130_fd_sc_hd__a211oi_1 _11709_ (.A1(\rbzero.floor_leak[5] ),
    .A2(_04810_),
    .B1(_04885_),
    .C1(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__clkbuf_4 _11710_ (.A(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__mux2_1 _11711_ (.A0(\rbzero.color_sky[0] ),
    .A1(\rbzero.color_floor[0] ),
    .S(_04825_),
    .X(_04901_));
 sky130_fd_sc_hd__buf_6 _11712_ (.A(_04812_),
    .X(_04902_));
 sky130_fd_sc_hd__buf_4 _11713_ (.A(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__buf_4 _11714_ (.A(_04891_),
    .X(_04904_));
 sky130_fd_sc_hd__clkbuf_4 _11715_ (.A(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__buf_4 _11716_ (.A(_04905_),
    .X(_04906_));
 sky130_fd_sc_hd__buf_4 _11717_ (.A(_04892_),
    .X(_04907_));
 sky130_fd_sc_hd__buf_6 _11718_ (.A(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__buf_6 _11719_ (.A(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__buf_6 _11720_ (.A(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__mux2_1 _11721_ (.A0(\rbzero.tex_r0[7] ),
    .A1(\rbzero.tex_r0[6] ),
    .S(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__buf_4 _11722_ (.A(_04827_),
    .X(_04912_));
 sky130_fd_sc_hd__buf_6 _11723_ (.A(_04892_),
    .X(_04913_));
 sky130_fd_sc_hd__clkbuf_8 _11724_ (.A(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__mux2_1 _11725_ (.A0(\rbzero.tex_r0[5] ),
    .A1(\rbzero.tex_r0[4] ),
    .S(_04914_),
    .X(_04915_));
 sky130_fd_sc_hd__or2_1 _11726_ (.A(_04912_),
    .B(_04915_),
    .X(_04916_));
 sky130_fd_sc_hd__nor3_4 _11727_ (.A(_04790_),
    .B(_04806_),
    .C(_04813_),
    .Y(_04917_));
 sky130_fd_sc_hd__buf_6 _11728_ (.A(_04917_),
    .X(_04918_));
 sky130_fd_sc_hd__clkbuf_8 _11729_ (.A(_04918_),
    .X(_04919_));
 sky130_fd_sc_hd__buf_4 _11730_ (.A(_04919_),
    .X(_04920_));
 sky130_fd_sc_hd__o211a_1 _11731_ (.A1(_04906_),
    .A2(_04911_),
    .B1(_04916_),
    .C1(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__buf_4 _11732_ (.A(_04827_),
    .X(_04922_));
 sky130_fd_sc_hd__buf_4 _11733_ (.A(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__buf_4 _11734_ (.A(_04914_),
    .X(_04924_));
 sky130_fd_sc_hd__mux2_1 _11735_ (.A0(\rbzero.tex_r0[1] ),
    .A1(\rbzero.tex_r0[0] ),
    .S(_04924_),
    .X(_04925_));
 sky130_fd_sc_hd__clkbuf_4 _11736_ (.A(_04785_),
    .X(_04926_));
 sky130_fd_sc_hd__buf_4 _11737_ (.A(_04926_),
    .X(_04927_));
 sky130_fd_sc_hd__clkbuf_4 _11738_ (.A(_04828_),
    .X(_04928_));
 sky130_fd_sc_hd__buf_4 _11739_ (.A(_04928_),
    .X(_04929_));
 sky130_fd_sc_hd__and3_1 _11740_ (.A(\rbzero.tex_r0[3] ),
    .B(_04927_),
    .C(_04929_),
    .X(_04930_));
 sky130_fd_sc_hd__buf_4 _11741_ (.A(_04893_),
    .X(_04931_));
 sky130_fd_sc_hd__buf_4 _11742_ (.A(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__buf_4 _11743_ (.A(_04932_),
    .X(_04933_));
 sky130_fd_sc_hd__buf_4 _11744_ (.A(_04891_),
    .X(_04934_));
 sky130_fd_sc_hd__buf_4 _11745_ (.A(_04934_),
    .X(_04935_));
 sky130_fd_sc_hd__a21o_1 _11746_ (.A1(\rbzero.tex_r0[2] ),
    .A2(_04933_),
    .B1(_04935_),
    .X(_04936_));
 sky130_fd_sc_hd__buf_6 _11747_ (.A(_04890_),
    .X(_04937_));
 sky130_fd_sc_hd__o221a_1 _11748_ (.A1(_04923_),
    .A2(_04925_),
    .B1(_04930_),
    .B2(_04936_),
    .C1(_04937_),
    .X(_04938_));
 sky130_fd_sc_hd__clkbuf_8 _11749_ (.A(_04814_),
    .X(_04939_));
 sky130_fd_sc_hd__buf_6 _11750_ (.A(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__buf_4 _11751_ (.A(_04940_),
    .X(_04941_));
 sky130_fd_sc_hd__mux2_1 _11752_ (.A0(\rbzero.tex_r0[9] ),
    .A1(\rbzero.tex_r0[8] ),
    .S(_04909_),
    .X(_04942_));
 sky130_fd_sc_hd__mux2_1 _11753_ (.A0(\rbzero.tex_r0[11] ),
    .A1(\rbzero.tex_r0[10] ),
    .S(_04909_),
    .X(_04943_));
 sky130_fd_sc_hd__buf_6 _11754_ (.A(_04827_),
    .X(_04944_));
 sky130_fd_sc_hd__mux2_1 _11755_ (.A0(_04942_),
    .A1(_04943_),
    .S(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__buf_4 _11756_ (.A(_04826_),
    .X(_04946_));
 sky130_fd_sc_hd__buf_6 _11757_ (.A(_04946_),
    .X(_04947_));
 sky130_fd_sc_hd__clkbuf_8 _11758_ (.A(_04908_),
    .X(_04948_));
 sky130_fd_sc_hd__mux2_1 _11759_ (.A0(\rbzero.tex_r0[13] ),
    .A1(\rbzero.tex_r0[12] ),
    .S(_04948_),
    .X(_04949_));
 sky130_fd_sc_hd__mux2_1 _11760_ (.A0(\rbzero.tex_r0[15] ),
    .A1(\rbzero.tex_r0[14] ),
    .S(_04908_),
    .X(_04950_));
 sky130_fd_sc_hd__or2_1 _11761_ (.A(_04934_),
    .B(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__clkbuf_8 _11762_ (.A(_04918_),
    .X(_04952_));
 sky130_fd_sc_hd__buf_6 _11763_ (.A(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__o211a_1 _11764_ (.A1(_04947_),
    .A2(_04949_),
    .B1(_04951_),
    .C1(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__buf_4 _11765_ (.A(_04889_),
    .X(_04955_));
 sky130_fd_sc_hd__a211o_1 _11766_ (.A1(_04941_),
    .A2(_04945_),
    .B1(_04954_),
    .C1(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__o311a_1 _11767_ (.A1(_04903_),
    .A2(_04921_),
    .A3(_04938_),
    .B1(_04956_),
    .C1(_04887_),
    .X(_04957_));
 sky130_fd_sc_hd__buf_6 _11768_ (.A(_04823_),
    .X(_04958_));
 sky130_fd_sc_hd__mux2_1 _11769_ (.A0(\rbzero.tex_r0[29] ),
    .A1(\rbzero.tex_r0[28] ),
    .S(_04914_),
    .X(_04959_));
 sky130_fd_sc_hd__mux2_1 _11770_ (.A0(\rbzero.tex_r0[31] ),
    .A1(\rbzero.tex_r0[30] ),
    .S(_04914_),
    .X(_04960_));
 sky130_fd_sc_hd__mux2_1 _11771_ (.A0(_04959_),
    .A1(_04960_),
    .S(_04944_),
    .X(_04961_));
 sky130_fd_sc_hd__mux2_1 _11772_ (.A0(\rbzero.tex_r0[25] ),
    .A1(\rbzero.tex_r0[24] ),
    .S(_04914_),
    .X(_04962_));
 sky130_fd_sc_hd__and3_1 _11773_ (.A(\rbzero.tex_r0[27] ),
    .B(_04927_),
    .C(_04929_),
    .X(_04963_));
 sky130_fd_sc_hd__clkbuf_8 _11774_ (.A(_04931_),
    .X(_04964_));
 sky130_fd_sc_hd__a21o_1 _11775_ (.A1(\rbzero.tex_r0[26] ),
    .A2(_04964_),
    .B1(_04934_),
    .X(_04965_));
 sky130_fd_sc_hd__o221a_1 _11776_ (.A1(_04912_),
    .A2(_04962_),
    .B1(_04963_),
    .B2(_04965_),
    .C1(_04940_),
    .X(_04966_));
 sky130_fd_sc_hd__buf_6 _11777_ (.A(_04889_),
    .X(_04967_));
 sky130_fd_sc_hd__a211o_1 _11778_ (.A1(_04920_),
    .A2(_04961_),
    .B1(_04966_),
    .C1(_04967_),
    .X(_04968_));
 sky130_fd_sc_hd__mux2_1 _11779_ (.A0(\rbzero.tex_r0[17] ),
    .A1(\rbzero.tex_r0[16] ),
    .S(_04914_),
    .X(_04969_));
 sky130_fd_sc_hd__mux2_1 _11780_ (.A0(\rbzero.tex_r0[19] ),
    .A1(\rbzero.tex_r0[18] ),
    .S(_04914_),
    .X(_04970_));
 sky130_fd_sc_hd__mux2_1 _11781_ (.A0(_04969_),
    .A1(_04970_),
    .S(_04944_),
    .X(_04971_));
 sky130_fd_sc_hd__mux2_1 _11782_ (.A0(\rbzero.tex_r0[21] ),
    .A1(\rbzero.tex_r0[20] ),
    .S(_04909_),
    .X(_04972_));
 sky130_fd_sc_hd__mux2_1 _11783_ (.A0(\rbzero.tex_r0[23] ),
    .A1(\rbzero.tex_r0[22] ),
    .S(_04913_),
    .X(_04973_));
 sky130_fd_sc_hd__or2_1 _11784_ (.A(_04934_),
    .B(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__o211a_1 _11785_ (.A1(_04947_),
    .A2(_04972_),
    .B1(_04974_),
    .C1(_04919_),
    .X(_04975_));
 sky130_fd_sc_hd__a211o_1 _11786_ (.A1(_04941_),
    .A2(_04971_),
    .B1(_04975_),
    .C1(_04902_),
    .X(_04976_));
 sky130_fd_sc_hd__a31o_1 _11787_ (.A1(_04958_),
    .A2(_04968_),
    .A3(_04976_),
    .B1(_04832_),
    .X(_04977_));
 sky130_fd_sc_hd__buf_6 _11788_ (.A(_04913_),
    .X(_04978_));
 sky130_fd_sc_hd__mux2_1 _11789_ (.A0(\rbzero.tex_r0[39] ),
    .A1(\rbzero.tex_r0[38] ),
    .S(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__mux2_1 _11790_ (.A0(\rbzero.tex_r0[37] ),
    .A1(\rbzero.tex_r0[36] ),
    .S(_04978_),
    .X(_04980_));
 sky130_fd_sc_hd__buf_4 _11791_ (.A(_04817_),
    .X(_04981_));
 sky130_fd_sc_hd__buf_4 _11792_ (.A(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__mux2_1 _11793_ (.A0(_04979_),
    .A1(_04980_),
    .S(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__mux2_1 _11794_ (.A0(\rbzero.tex_r0[33] ),
    .A1(\rbzero.tex_r0[32] ),
    .S(_04978_),
    .X(_04984_));
 sky130_fd_sc_hd__mux2_1 _11795_ (.A0(\rbzero.tex_r0[35] ),
    .A1(\rbzero.tex_r0[34] ),
    .S(_04978_),
    .X(_04985_));
 sky130_fd_sc_hd__mux2_1 _11796_ (.A0(_04984_),
    .A1(_04985_),
    .S(_04922_),
    .X(_04986_));
 sky130_fd_sc_hd__mux2_1 _11797_ (.A0(_04983_),
    .A1(_04986_),
    .S(_04937_),
    .X(_04987_));
 sky130_fd_sc_hd__mux2_1 _11798_ (.A0(\rbzero.tex_r0[47] ),
    .A1(\rbzero.tex_r0[46] ),
    .S(_04910_),
    .X(_04988_));
 sky130_fd_sc_hd__mux2_1 _11799_ (.A0(\rbzero.tex_r0[45] ),
    .A1(\rbzero.tex_r0[44] ),
    .S(_04948_),
    .X(_04989_));
 sky130_fd_sc_hd__or2_1 _11800_ (.A(_04947_),
    .B(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__o211a_1 _11801_ (.A1(_04906_),
    .A2(_04988_),
    .B1(_04990_),
    .C1(_04920_),
    .X(_04991_));
 sky130_fd_sc_hd__mux2_1 _11802_ (.A0(\rbzero.tex_r0[41] ),
    .A1(\rbzero.tex_r0[40] ),
    .S(_04948_),
    .X(_04992_));
 sky130_fd_sc_hd__mux2_1 _11803_ (.A0(\rbzero.tex_r0[43] ),
    .A1(\rbzero.tex_r0[42] ),
    .S(_04948_),
    .X(_04993_));
 sky130_fd_sc_hd__mux2_1 _11804_ (.A0(_04992_),
    .A1(_04993_),
    .S(_04912_),
    .X(_04994_));
 sky130_fd_sc_hd__a21o_1 _11805_ (.A1(_04941_),
    .A2(_04994_),
    .B1(_04955_),
    .X(_04995_));
 sky130_fd_sc_hd__o221a_1 _11806_ (.A1(_04903_),
    .A2(_04987_),
    .B1(_04991_),
    .B2(_04995_),
    .C1(_04887_),
    .X(_04996_));
 sky130_fd_sc_hd__mux2_1 _11807_ (.A0(\rbzero.tex_r0[53] ),
    .A1(\rbzero.tex_r0[52] ),
    .S(_04909_),
    .X(_04997_));
 sky130_fd_sc_hd__mux2_1 _11808_ (.A0(\rbzero.tex_r0[55] ),
    .A1(\rbzero.tex_r0[54] ),
    .S(_04909_),
    .X(_04998_));
 sky130_fd_sc_hd__mux2_1 _11809_ (.A0(_04997_),
    .A1(_04998_),
    .S(_04944_),
    .X(_04999_));
 sky130_fd_sc_hd__mux2_1 _11810_ (.A0(\rbzero.tex_r0[49] ),
    .A1(\rbzero.tex_r0[48] ),
    .S(_04914_),
    .X(_05000_));
 sky130_fd_sc_hd__and3_1 _11811_ (.A(\rbzero.tex_r0[51] ),
    .B(_04927_),
    .C(_04929_),
    .X(_05001_));
 sky130_fd_sc_hd__buf_4 _11812_ (.A(_04978_),
    .X(_05002_));
 sky130_fd_sc_hd__a21o_1 _11813_ (.A1(\rbzero.tex_r0[50] ),
    .A2(_05002_),
    .B1(_04934_),
    .X(_05003_));
 sky130_fd_sc_hd__o221a_1 _11814_ (.A1(_04912_),
    .A2(_05000_),
    .B1(_05001_),
    .B2(_05003_),
    .C1(_04940_),
    .X(_05004_));
 sky130_fd_sc_hd__a211o_1 _11815_ (.A1(_04920_),
    .A2(_04999_),
    .B1(_05004_),
    .C1(_04902_),
    .X(_05005_));
 sky130_fd_sc_hd__mux2_1 _11816_ (.A0(\rbzero.tex_r0[57] ),
    .A1(\rbzero.tex_r0[56] ),
    .S(_04909_),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_1 _11817_ (.A0(\rbzero.tex_r0[59] ),
    .A1(\rbzero.tex_r0[58] ),
    .S(_04909_),
    .X(_05007_));
 sky130_fd_sc_hd__mux2_1 _11818_ (.A0(_05006_),
    .A1(_05007_),
    .S(_04944_),
    .X(_05008_));
 sky130_fd_sc_hd__buf_4 _11819_ (.A(_04907_),
    .X(_05009_));
 sky130_fd_sc_hd__buf_6 _11820_ (.A(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__and2_1 _11821_ (.A(\rbzero.tex_r0[62] ),
    .B(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__a31o_1 _11822_ (.A1(\rbzero.tex_r0[63] ),
    .A2(_04927_),
    .A3(_04929_),
    .B1(_04904_),
    .X(_05012_));
 sky130_fd_sc_hd__mux2_1 _11823_ (.A0(\rbzero.tex_r0[61] ),
    .A1(\rbzero.tex_r0[60] ),
    .S(_04909_),
    .X(_05013_));
 sky130_fd_sc_hd__o221a_1 _11824_ (.A1(_05011_),
    .A2(_05012_),
    .B1(_05013_),
    .B2(_04947_),
    .C1(_04919_),
    .X(_05014_));
 sky130_fd_sc_hd__a211o_1 _11825_ (.A1(_04941_),
    .A2(_05008_),
    .B1(_05014_),
    .C1(_04955_),
    .X(_05015_));
 sky130_fd_sc_hd__a31o_1 _11826_ (.A1(_04958_),
    .A2(_05005_),
    .A3(_05015_),
    .B1(_04810_),
    .X(_05016_));
 sky130_fd_sc_hd__clkinv_4 _11827_ (.A(net42),
    .Y(_05017_));
 sky130_fd_sc_hd__o221a_2 _11828_ (.A1(_04957_),
    .A2(_04977_),
    .B1(_04996_),
    .B2(_05016_),
    .C1(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__or2b_1 _11829_ (.A(\rbzero.row_render.wall[1] ),
    .B_N(\rbzero.row_render.wall[0] ),
    .X(_05019_));
 sky130_fd_sc_hd__or2b_1 _11830_ (.A(\rbzero.row_render.wall[0] ),
    .B_N(\rbzero.row_render.wall[1] ),
    .X(_05020_));
 sky130_fd_sc_hd__inv_2 _11831_ (.A(\rbzero.row_render.texu[3] ),
    .Y(_05021_));
 sky130_fd_sc_hd__nand2_1 _11832_ (.A(\rbzero.row_render.texu[2] ),
    .B(\rbzero.row_render.texu[1] ),
    .Y(_05022_));
 sky130_fd_sc_hd__o21ai_1 _11833_ (.A1(_05021_),
    .A2(_05022_),
    .B1(_04819_),
    .Y(_05023_));
 sky130_fd_sc_hd__nor2_1 _11834_ (.A(\rbzero.row_render.texu[2] ),
    .B(\rbzero.row_render.texu[1] ),
    .Y(_05024_));
 sky130_fd_sc_hd__a32o_1 _11835_ (.A1(_04812_),
    .A2(_04917_),
    .A3(_04826_),
    .B1(_05024_),
    .B2(_05021_),
    .X(_05025_));
 sky130_fd_sc_hd__inv_2 _11836_ (.A(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__inv_2 _11837_ (.A(\rbzero.row_render.side ),
    .Y(_05027_));
 sky130_fd_sc_hd__a41o_1 _11838_ (.A1(\rbzero.row_render.wall[0] ),
    .A2(\rbzero.row_render.wall[1] ),
    .A3(_05023_),
    .A4(_05026_),
    .B1(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__and3_1 _11839_ (.A(_05027_),
    .B(\rbzero.row_render.wall[0] ),
    .C(_05026_),
    .X(_05029_));
 sky130_fd_sc_hd__nand3_1 _11840_ (.A(\rbzero.row_render.wall[1] ),
    .B(_05023_),
    .C(_05029_),
    .Y(_05030_));
 sky130_fd_sc_hd__clkbuf_4 _11841_ (.A(_04829_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_4 _11842_ (.A(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__or3b_1 _11843_ (.A(_05032_),
    .B(_04818_),
    .C_N(\rbzero.row_render.texu[0] ),
    .X(_05033_));
 sky130_fd_sc_hd__o31a_1 _11844_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(\rbzero.row_render.texu[3] ),
    .A3(_05022_),
    .B1(_04889_),
    .X(_05034_));
 sky130_fd_sc_hd__a31o_1 _11845_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(\rbzero.row_render.texu[3] ),
    .A3(_05024_),
    .B1(_04889_),
    .X(_05035_));
 sky130_fd_sc_hd__or3b_1 _11846_ (.A(\rbzero.row_render.texu[0] ),
    .B(_05034_),
    .C_N(_05035_),
    .X(_05036_));
 sky130_fd_sc_hd__o31ai_2 _11847_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_04818_),
    .A3(_05031_),
    .B1(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__nor2_1 _11848_ (.A(\rbzero.row_render.side ),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__a21oi_1 _11849_ (.A1(\rbzero.row_render.side ),
    .A2(_05033_),
    .B1(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__nor2_1 _11850_ (.A(_05020_),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__a31o_1 _11851_ (.A1(_05020_),
    .A2(_05028_),
    .A3(_05030_),
    .B1(_05040_),
    .X(_05041_));
 sky130_fd_sc_hd__and2b_1 _11852_ (.A_N(\rbzero.row_render.wall[1] ),
    .B(\rbzero.row_render.wall[0] ),
    .X(_05042_));
 sky130_fd_sc_hd__a21o_1 _11853_ (.A1(_05027_),
    .A2(_05042_),
    .B1(_05017_),
    .X(_05043_));
 sky130_fd_sc_hd__a21o_1 _11854_ (.A1(_05019_),
    .A2(_05041_),
    .B1(_05043_),
    .X(_05044_));
 sky130_fd_sc_hd__nand2_1 _11855_ (.A(_04900_),
    .B(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__o22a_1 _11856_ (.A1(_04900_),
    .A2(_04901_),
    .B1(_05018_),
    .B2(_05045_),
    .X(_05046_));
 sky130_fd_sc_hd__nor3_2 _11857_ (.A(_04696_),
    .B(_04697_),
    .C(_04701_),
    .Y(_05047_));
 sky130_fd_sc_hd__o22a_1 _11858_ (.A1(_04703_),
    .A2(_04745_),
    .B1(_05046_),
    .B2(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__nor2_1 _11859_ (.A(_04650_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__and3_4 _11860_ (.A(\rbzero.trace_state[3] ),
    .B(_04429_),
    .C(_04436_),
    .X(_05050_));
 sky130_fd_sc_hd__a21o_1 _11861_ (.A1(\rbzero.trace_state[0] ),
    .A2(_05050_),
    .B1(_04635_),
    .X(_05051_));
 sky130_fd_sc_hd__o21ai_1 _11862_ (.A1(_04661_),
    .A2(_05049_),
    .B1(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__o21a_4 _11863_ (.A1(\gpout0.hpos[7] ),
    .A2(\gpout0.hpos[8] ),
    .B1(\gpout0.hpos[9] ),
    .X(_05053_));
 sky130_fd_sc_hd__and3_1 _11864_ (.A(\gpout0.vpos[7] ),
    .B(_04648_),
    .C(_04656_),
    .X(_05054_));
 sky130_fd_sc_hd__a21o_4 _11865_ (.A1(\gpout0.vpos[8] ),
    .A2(_05054_),
    .B1(\gpout0.vpos[9] ),
    .X(_05055_));
 sky130_fd_sc_hd__nor2_2 _11866_ (.A(_05053_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__o211a_4 _11867_ (.A1(\rbzero.trace_state[0] ),
    .A2(_04635_),
    .B1(_05052_),
    .C1(_05056_),
    .X(_05057_));
 sky130_fd_sc_hd__buf_6 _11868_ (.A(net45),
    .X(_05058_));
 sky130_fd_sc_hd__mux2_2 _11869_ (.A0(\reg_rgb[6] ),
    .A1(_05057_),
    .S(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__clkbuf_1 _11870_ (.A(_05059_),
    .X(net68));
 sky130_fd_sc_hd__nor2_1 _11871_ (.A(_04412_),
    .B(_04636_),
    .Y(_05060_));
 sky130_fd_sc_hd__or2_2 _11872_ (.A(_04637_),
    .B(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__nor2_1 _11873_ (.A(_04415_),
    .B(_04632_),
    .Y(_05062_));
 sky130_fd_sc_hd__or4bb_1 _11874_ (.A(_04824_),
    .B(_05062_),
    .C_N(_04424_),
    .D_N(_03977_),
    .X(_05063_));
 sky130_fd_sc_hd__nor2_2 _11875_ (.A(_04656_),
    .B(_04655_),
    .Y(_05064_));
 sky130_fd_sc_hd__nor2_1 _11876_ (.A(\gpout0.hpos[7] ),
    .B(_04639_),
    .Y(_05065_));
 sky130_fd_sc_hd__or2_1 _11877_ (.A(_04640_),
    .B(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__nor2_1 _11878_ (.A(\gpout0.hpos[4] ),
    .B(_05061_),
    .Y(_05067_));
 sky130_fd_sc_hd__o21ba_1 _11879_ (.A1(_04638_),
    .A2(_04699_),
    .B1_N(_04639_),
    .X(_05068_));
 sky130_fd_sc_hd__mux2_1 _11880_ (.A0(\gpout0.hpos[6] ),
    .A1(_04630_),
    .S(_04636_),
    .X(_05069_));
 sky130_fd_sc_hd__or3_1 _11881_ (.A(_05067_),
    .B(_05068_),
    .C(_05069_),
    .X(_05070_));
 sky130_fd_sc_hd__a2bb2o_1 _11882_ (.A1_N(_05067_),
    .A2_N(_05068_),
    .B1(\gpout0.hpos[6] ),
    .B2(\gpout0.hpos[5] ),
    .X(_05071_));
 sky130_fd_sc_hd__nand2_1 _11883_ (.A(_05070_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__xor2_2 _11884_ (.A(_05066_),
    .B(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__nor2_1 _11885_ (.A(_04421_),
    .B(_04636_),
    .Y(_05074_));
 sky130_fd_sc_hd__a21oi_4 _11886_ (.A1(_04424_),
    .A2(_04636_),
    .B1(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__or2_1 _11887_ (.A(_05066_),
    .B(_05070_),
    .X(_05076_));
 sky130_fd_sc_hd__or3b_1 _11888_ (.A(_04641_),
    .B(_05053_),
    .C_N(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__or2b_1 _11889_ (.A(_05077_),
    .B_N(_05061_),
    .X(_05078_));
 sky130_fd_sc_hd__nand2_1 _11890_ (.A(_04415_),
    .B(_04636_),
    .Y(_05079_));
 sky130_fd_sc_hd__nand3b_4 _11891_ (.A_N(_05078_),
    .B(_05079_),
    .C(_04638_),
    .Y(_05080_));
 sky130_fd_sc_hd__a21oi_1 _11892_ (.A1(_04638_),
    .A2(_05079_),
    .B1(_05078_),
    .Y(_05081_));
 sky130_fd_sc_hd__or2b_2 _11893_ (.A(_05075_),
    .B_N(_05081_),
    .X(_05082_));
 sky130_fd_sc_hd__or2_1 _11894_ (.A(_05061_),
    .B(_05077_),
    .X(_05083_));
 sky130_fd_sc_hd__inv_2 _11895_ (.A(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__nand3_2 _11896_ (.A(_04578_),
    .B(_05075_),
    .C(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__or3_2 _11897_ (.A(\gpout0.hpos[4] ),
    .B(_05075_),
    .C(_05083_),
    .X(_05086_));
 sky130_fd_sc_hd__o21bai_1 _11898_ (.A1(_05066_),
    .A2(_05071_),
    .B1_N(_04640_),
    .Y(_05087_));
 sky130_fd_sc_hd__xor2_1 _11899_ (.A(\gpout0.hpos[8] ),
    .B(_05087_),
    .X(_05088_));
 sky130_fd_sc_hd__or2b_2 _11900_ (.A(_05088_),
    .B_N(_05069_),
    .X(_05089_));
 sky130_fd_sc_hd__a41o_1 _11901_ (.A1(_05080_),
    .A2(_05082_),
    .A3(_05085_),
    .A4(_05086_),
    .B1(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__o21ai_1 _11902_ (.A1(_05075_),
    .A2(_05080_),
    .B1(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__o21bai_1 _11903_ (.A1(_05076_),
    .A2(_05088_),
    .B1_N(_05069_),
    .Y(_05092_));
 sky130_fd_sc_hd__a21o_4 _11904_ (.A1(_05076_),
    .A2(_05088_),
    .B1(_05092_),
    .X(_05093_));
 sky130_fd_sc_hd__nand2_1 _11905_ (.A(_05075_),
    .B(_05081_),
    .Y(_05094_));
 sky130_fd_sc_hd__nor2_1 _11906_ (.A(_05093_),
    .B(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__nor2_1 _11907_ (.A(_05085_),
    .B(_05093_),
    .Y(_05096_));
 sky130_fd_sc_hd__or3b_2 _11908_ (.A(_05083_),
    .B(\gpout0.hpos[4] ),
    .C_N(_05075_),
    .X(_05097_));
 sky130_fd_sc_hd__nor2_1 _11909_ (.A(_05093_),
    .B(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__or3_1 _11910_ (.A(_05095_),
    .B(_05096_),
    .C(_05098_),
    .X(_05099_));
 sky130_fd_sc_hd__nor3_1 _11911_ (.A(_04414_),
    .B(_05075_),
    .C(_05083_),
    .Y(_05100_));
 sky130_fd_sc_hd__and2_1 _11912_ (.A(_05073_),
    .B(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__or2_1 _11913_ (.A(_04411_),
    .B(_05080_),
    .X(_05102_));
 sky130_fd_sc_hd__nor2_1 _11914_ (.A(_05093_),
    .B(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__or3_1 _11915_ (.A(_05099_),
    .B(_05101_),
    .C(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__a21o_2 _11916_ (.A1(_05073_),
    .A2(_05091_),
    .B1(_05104_),
    .X(_05105_));
 sky130_fd_sc_hd__clkbuf_4 _11917_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .X(_05106_));
 sky130_fd_sc_hd__nor3_4 _11918_ (.A(_05075_),
    .B(_05080_),
    .C(_05093_),
    .Y(_05107_));
 sky130_fd_sc_hd__nor2_4 _11919_ (.A(_05086_),
    .B(_05093_),
    .Y(_05108_));
 sky130_fd_sc_hd__a22o_1 _11920_ (.A1(_05106_),
    .A2(_05107_),
    .B1(_05108_),
    .B2(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(_05109_));
 sky130_fd_sc_hd__and2b_2 _11921_ (.A_N(_05093_),
    .B(_05100_),
    .X(_05110_));
 sky130_fd_sc_hd__buf_4 _11922_ (.A(\rbzero.debug_overlay.vplaneX[-5] ),
    .X(_05111_));
 sky130_fd_sc_hd__nor2_4 _11923_ (.A(_05089_),
    .B(_05097_),
    .Y(_05112_));
 sky130_fd_sc_hd__nor2_4 _11924_ (.A(_05089_),
    .B(_05094_),
    .Y(_05113_));
 sky130_fd_sc_hd__a221o_1 _11925_ (.A1(_05111_),
    .A2(_05112_),
    .B1(_05113_),
    .B2(\rbzero.debug_overlay.vplaneX[-4] ),
    .C1(_04652_),
    .X(_05114_));
 sky130_fd_sc_hd__nor2_4 _11926_ (.A(_05082_),
    .B(_05093_),
    .Y(_05115_));
 sky130_fd_sc_hd__or2_4 _11927_ (.A(_05073_),
    .B(_05089_),
    .X(_05116_));
 sky130_fd_sc_hd__nor2_4 _11928_ (.A(_05082_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__nor2_4 _11929_ (.A(_05085_),
    .B(_05116_),
    .Y(_05118_));
 sky130_fd_sc_hd__a22o_1 _11930_ (.A1(\rbzero.debug_overlay.vplaneX[-8] ),
    .A2(_05117_),
    .B1(_05118_),
    .B2(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(_05119_));
 sky130_fd_sc_hd__clkbuf_4 _11931_ (.A(\rbzero.debug_overlay.vplaneX[-6] ),
    .X(_05120_));
 sky130_fd_sc_hd__nor2_4 _11932_ (.A(_05102_),
    .B(_05116_),
    .Y(_05121_));
 sky130_fd_sc_hd__nor2_4 _11933_ (.A(_05086_),
    .B(_05116_),
    .Y(_05122_));
 sky130_fd_sc_hd__a22o_1 _11934_ (.A1(_05120_),
    .A2(_05121_),
    .B1(_05122_),
    .B2(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_05123_));
 sky130_fd_sc_hd__a211o_1 _11935_ (.A1(\rbzero.debug_overlay.vplaneX[0] ),
    .A2(_05115_),
    .B1(_05119_),
    .C1(_05123_),
    .X(_05124_));
 sky130_fd_sc_hd__a211o_1 _11936_ (.A1(\rbzero.debug_overlay.vplaneX[-3] ),
    .A2(_05110_),
    .B1(_05114_),
    .C1(_05124_),
    .X(_05125_));
 sky130_fd_sc_hd__a211o_2 _11937_ (.A1(\rbzero.debug_overlay.vplaneX[10] ),
    .A2(_05105_),
    .B1(_05109_),
    .C1(_05125_),
    .X(_05126_));
 sky130_fd_sc_hd__buf_2 _11938_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .X(_05127_));
 sky130_fd_sc_hd__a22o_1 _11939_ (.A1(\rbzero.debug_overlay.vplaneY[-1] ),
    .A2(_05108_),
    .B1(_05115_),
    .B2(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_05128_));
 sky130_fd_sc_hd__clkbuf_4 _11940_ (.A(\rbzero.debug_overlay.vplaneY[-6] ),
    .X(_05129_));
 sky130_fd_sc_hd__a22o_1 _11941_ (.A1(_05129_),
    .A2(_05121_),
    .B1(_05122_),
    .B2(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_05130_));
 sky130_fd_sc_hd__a221o_1 _11942_ (.A1(\rbzero.debug_overlay.vplaneY[-8] ),
    .A2(_05117_),
    .B1(_05118_),
    .B2(\rbzero.debug_overlay.vplaneY[-7] ),
    .C1(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__buf_2 _11943_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .X(_05132_));
 sky130_fd_sc_hd__a21bo_1 _11944_ (.A1(\rbzero.debug_overlay.vplaneY[-5] ),
    .A2(_05112_),
    .B1_N(_04652_),
    .X(_05133_));
 sky130_fd_sc_hd__a221o_1 _11945_ (.A1(\rbzero.debug_overlay.vplaneY[-2] ),
    .A2(_05107_),
    .B1(_05113_),
    .B2(_05132_),
    .C1(_05133_),
    .X(_05134_));
 sky130_fd_sc_hd__a2111o_1 _11946_ (.A1(\rbzero.debug_overlay.vplaneY[-3] ),
    .A2(_05110_),
    .B1(_05128_),
    .C1(_05131_),
    .D1(_05134_),
    .X(_05135_));
 sky130_fd_sc_hd__a21o_2 _11947_ (.A1(_05127_),
    .A2(_05105_),
    .B1(_05135_),
    .X(_05136_));
 sky130_fd_sc_hd__a22o_1 _11948_ (.A1(\rbzero.debug_overlay.facingY[-3] ),
    .A2(_05110_),
    .B1(_05108_),
    .B2(\rbzero.debug_overlay.facingY[-1] ),
    .X(_05137_));
 sky130_fd_sc_hd__a22o_1 _11949_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_05121_),
    .B1(_05118_),
    .B2(\rbzero.debug_overlay.facingY[-7] ),
    .X(_05138_));
 sky130_fd_sc_hd__a22o_1 _11950_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_05112_),
    .B1(_05113_),
    .B2(\rbzero.debug_overlay.facingY[-4] ),
    .X(_05139_));
 sky130_fd_sc_hd__a221o_1 _11951_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(_05107_),
    .B1(_05122_),
    .B2(\rbzero.debug_overlay.facingY[-9] ),
    .C1(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__a211o_1 _11952_ (.A1(\rbzero.debug_overlay.facingY[-8] ),
    .A2(_05117_),
    .B1(_05138_),
    .C1(_05140_),
    .X(_05141_));
 sky130_fd_sc_hd__a211o_1 _11953_ (.A1(\rbzero.debug_overlay.facingY[0] ),
    .A2(_05115_),
    .B1(_05137_),
    .C1(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__a21oi_2 _11954_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(_05105_),
    .B1(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__nor3_1 _11955_ (.A(_04731_),
    .B(_04654_),
    .C(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__a41o_1 _11956_ (.A1(_04657_),
    .A2(_04651_),
    .A3(_05126_),
    .A4(_05136_),
    .B1(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__a22o_1 _11957_ (.A1(\rbzero.debug_overlay.facingX[-8] ),
    .A2(_05117_),
    .B1(_05122_),
    .B2(\rbzero.debug_overlay.facingX[-9] ),
    .X(_05146_));
 sky130_fd_sc_hd__a22o_1 _11958_ (.A1(\rbzero.debug_overlay.facingX[-6] ),
    .A2(_05121_),
    .B1(_05118_),
    .B2(\rbzero.debug_overlay.facingX[-7] ),
    .X(_05147_));
 sky130_fd_sc_hd__or2_1 _11959_ (.A(_05146_),
    .B(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__a21bo_1 _11960_ (.A1(\rbzero.debug_overlay.facingX[-5] ),
    .A2(_05112_),
    .B1_N(_05064_),
    .X(_05149_));
 sky130_fd_sc_hd__a221o_1 _11961_ (.A1(\rbzero.debug_overlay.facingX[-2] ),
    .A2(_05107_),
    .B1(_05113_),
    .B2(\rbzero.debug_overlay.facingX[-4] ),
    .C1(_05149_),
    .X(_05150_));
 sky130_fd_sc_hd__a22o_1 _11962_ (.A1(\rbzero.debug_overlay.facingX[-3] ),
    .A2(_05110_),
    .B1(_05108_),
    .B2(\rbzero.debug_overlay.facingX[-1] ),
    .X(_05151_));
 sky130_fd_sc_hd__a221o_1 _11963_ (.A1(\rbzero.debug_overlay.facingX[10] ),
    .A2(_05105_),
    .B1(_05115_),
    .B2(\rbzero.debug_overlay.facingX[0] ),
    .C1(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__or3_2 _11964_ (.A(_05148_),
    .B(_05150_),
    .C(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__o21ai_1 _11965_ (.A1(_05064_),
    .A2(_05145_),
    .B1(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__a22o_1 _11966_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_05098_),
    .B1(_05115_),
    .B2(\rbzero.debug_overlay.playerX[0] ),
    .X(_05155_));
 sky130_fd_sc_hd__a22o_1 _11967_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_05096_),
    .B1(_05110_),
    .B2(\rbzero.debug_overlay.playerX[-3] ),
    .X(_05156_));
 sky130_fd_sc_hd__a221o_1 _11968_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_05095_),
    .B1(_05108_),
    .B2(\rbzero.debug_overlay.playerX[-1] ),
    .C1(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__a22o_1 _11969_ (.A1(\rbzero.debug_overlay.playerX[-6] ),
    .A2(_05121_),
    .B1(_05118_),
    .B2(\rbzero.debug_overlay.playerX[-7] ),
    .X(_05158_));
 sky130_fd_sc_hd__a221o_1 _11970_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(_05117_),
    .B1(_05122_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__a221o_1 _11971_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(_05101_),
    .B1(_05112_),
    .B2(\rbzero.debug_overlay.playerX[-5] ),
    .C1(_04646_),
    .X(_05160_));
 sky130_fd_sc_hd__a221o_1 _11972_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_05107_),
    .B1(_05113_),
    .B2(\rbzero.debug_overlay.playerX[-4] ),
    .C1(_05160_),
    .X(_05161_));
 sky130_fd_sc_hd__or3_1 _11973_ (.A(_05157_),
    .B(_05159_),
    .C(_05161_),
    .X(_05162_));
 sky130_fd_sc_hd__a211oi_1 _11974_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_05103_),
    .B1(_05155_),
    .C1(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__a22o_1 _11975_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_05103_),
    .B1(_05115_),
    .B2(\rbzero.debug_overlay.playerY[0] ),
    .X(_05164_));
 sky130_fd_sc_hd__a22o_1 _11976_ (.A1(\rbzero.debug_overlay.playerY[-6] ),
    .A2(_05121_),
    .B1(_05117_),
    .B2(\rbzero.debug_overlay.playerY[-8] ),
    .X(_05165_));
 sky130_fd_sc_hd__a22o_1 _11977_ (.A1(\rbzero.debug_overlay.playerY[-9] ),
    .A2(_05122_),
    .B1(_05118_),
    .B2(\rbzero.debug_overlay.playerY[-7] ),
    .X(_05166_));
 sky130_fd_sc_hd__a22o_1 _11978_ (.A1(\rbzero.debug_overlay.playerY[4] ),
    .A2(_05095_),
    .B1(_05096_),
    .B2(\rbzero.debug_overlay.playerY[1] ),
    .X(_05167_));
 sky130_fd_sc_hd__a221o_1 _11979_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_05107_),
    .B1(_05110_),
    .B2(\rbzero.debug_overlay.playerY[-3] ),
    .C1(_05167_),
    .X(_05168_));
 sky130_fd_sc_hd__or3b_1 _11980_ (.A(_04656_),
    .B(\gpout0.vpos[4] ),
    .C_N(\gpout0.vpos[3] ),
    .X(_05169_));
 sky130_fd_sc_hd__a221o_1 _11981_ (.A1(\rbzero.debug_overlay.playerY[5] ),
    .A2(_05101_),
    .B1(_05113_),
    .B2(\rbzero.debug_overlay.playerY[-4] ),
    .C1(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__a221o_1 _11982_ (.A1(\rbzero.debug_overlay.playerY[-1] ),
    .A2(_05108_),
    .B1(_05112_),
    .B2(\rbzero.debug_overlay.playerY[-5] ),
    .C1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__or4_1 _11983_ (.A(_05165_),
    .B(_05166_),
    .C(_05168_),
    .D(_05171_),
    .X(_05172_));
 sky130_fd_sc_hd__a211o_1 _11984_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_05098_),
    .B1(_05164_),
    .C1(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__or3b_1 _11985_ (.A(_04659_),
    .B(_05163_),
    .C_N(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__a21o_1 _11986_ (.A1(_04645_),
    .A2(_05154_),
    .B1(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__o311a_1 _11987_ (.A1(_04589_),
    .A2(_05061_),
    .A3(_05063_),
    .B1(_05175_),
    .C1(_04650_),
    .X(_05176_));
 sky130_fd_sc_hd__a21o_1 _11988_ (.A1(\rbzero.row_render.side ),
    .A2(_05037_),
    .B1(_05020_),
    .X(_05177_));
 sky130_fd_sc_hd__o21ai_1 _11989_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_04958_),
    .B1(_05042_),
    .Y(_05178_));
 sky130_fd_sc_hd__a21oi_1 _11990_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_04958_),
    .B1(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__a31o_1 _11991_ (.A1(_05019_),
    .A2(_05030_),
    .A3(_05177_),
    .B1(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__clkbuf_4 _11992_ (.A(_04910_),
    .X(_05181_));
 sky130_fd_sc_hd__buf_4 _11993_ (.A(_04830_),
    .X(_05182_));
 sky130_fd_sc_hd__or2_1 _11994_ (.A(\rbzero.tex_r1[14] ),
    .B(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__o211a_1 _11995_ (.A1(\rbzero.tex_r1[15] ),
    .A2(_04933_),
    .B1(_05183_),
    .C1(_04923_),
    .X(_05184_));
 sky130_fd_sc_hd__buf_4 _11996_ (.A(_04982_),
    .X(_05185_));
 sky130_fd_sc_hd__buf_4 _11997_ (.A(_04831_),
    .X(_05186_));
 sky130_fd_sc_hd__a31o_1 _11998_ (.A1(\rbzero.tex_r1[13] ),
    .A2(_05185_),
    .A3(_05186_),
    .B1(_04937_),
    .X(_05187_));
 sky130_fd_sc_hd__a311o_1 _11999_ (.A1(\rbzero.tex_r1[12] ),
    .A2(_04906_),
    .A3(_05181_),
    .B1(_05184_),
    .C1(_05187_),
    .X(_05188_));
 sky130_fd_sc_hd__or2_1 _12000_ (.A(\rbzero.tex_r1[10] ),
    .B(_05182_),
    .X(_05189_));
 sky130_fd_sc_hd__buf_4 _12001_ (.A(_04826_),
    .X(_05190_));
 sky130_fd_sc_hd__buf_4 _12002_ (.A(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__o211a_1 _12003_ (.A1(\rbzero.tex_r1[11] ),
    .A2(_04933_),
    .B1(_05189_),
    .C1(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__a31o_1 _12004_ (.A1(\rbzero.tex_r1[9] ),
    .A2(_05185_),
    .A3(_05186_),
    .B1(_04953_),
    .X(_05193_));
 sky130_fd_sc_hd__a311o_1 _12005_ (.A1(\rbzero.tex_r1[8] ),
    .A2(_04906_),
    .A3(_05181_),
    .B1(_05192_),
    .C1(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__clkbuf_4 _12006_ (.A(_04924_),
    .X(_05195_));
 sky130_fd_sc_hd__or2_1 _12007_ (.A(\rbzero.tex_r1[6] ),
    .B(_05182_),
    .X(_05196_));
 sky130_fd_sc_hd__o211a_1 _12008_ (.A1(\rbzero.tex_r1[7] ),
    .A2(_05195_),
    .B1(_05196_),
    .C1(_04923_),
    .X(_05197_));
 sky130_fd_sc_hd__buf_4 _12009_ (.A(_04817_),
    .X(_05198_));
 sky130_fd_sc_hd__buf_4 _12010_ (.A(_05198_),
    .X(_05199_));
 sky130_fd_sc_hd__a31o_1 _12011_ (.A1(\rbzero.tex_r1[5] ),
    .A2(_05199_),
    .A3(_05032_),
    .B1(_04890_),
    .X(_05200_));
 sky130_fd_sc_hd__a31o_1 _12012_ (.A1(\rbzero.tex_r1[4] ),
    .A2(_05185_),
    .A3(_05195_),
    .B1(_05200_),
    .X(_05201_));
 sky130_fd_sc_hd__or2_1 _12013_ (.A(\rbzero.tex_r1[2] ),
    .B(_05032_),
    .X(_05202_));
 sky130_fd_sc_hd__o211a_1 _12014_ (.A1(\rbzero.tex_r1[3] ),
    .A2(_05195_),
    .B1(_05202_),
    .C1(_04923_),
    .X(_05203_));
 sky130_fd_sc_hd__a31o_1 _12015_ (.A1(\rbzero.tex_r1[1] ),
    .A2(_04982_),
    .A3(_05032_),
    .B1(_04919_),
    .X(_05204_));
 sky130_fd_sc_hd__a31o_1 _12016_ (.A1(\rbzero.tex_r1[0] ),
    .A2(_05185_),
    .A3(_05181_),
    .B1(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__o221a_1 _12017_ (.A1(_05197_),
    .A2(_05201_),
    .B1(_05203_),
    .B2(_05205_),
    .C1(_04955_),
    .X(_05206_));
 sky130_fd_sc_hd__a311o_1 _12018_ (.A1(_04903_),
    .A2(_05188_),
    .A3(_05194_),
    .B1(_04958_),
    .C1(_05206_),
    .X(_05207_));
 sky130_fd_sc_hd__or2_1 _12019_ (.A(\rbzero.tex_r1[22] ),
    .B(_05182_),
    .X(_05208_));
 sky130_fd_sc_hd__o211a_1 _12020_ (.A1(\rbzero.tex_r1[23] ),
    .A2(_04933_),
    .B1(_05208_),
    .C1(_04923_),
    .X(_05209_));
 sky130_fd_sc_hd__a31o_1 _12021_ (.A1(\rbzero.tex_r1[21] ),
    .A2(_05185_),
    .A3(_05186_),
    .B1(_04937_),
    .X(_05210_));
 sky130_fd_sc_hd__a311o_1 _12022_ (.A1(\rbzero.tex_r1[20] ),
    .A2(_04906_),
    .A3(_05181_),
    .B1(_05209_),
    .C1(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__or2_1 _12023_ (.A(\rbzero.tex_r1[18] ),
    .B(_05182_),
    .X(_05212_));
 sky130_fd_sc_hd__o211a_1 _12024_ (.A1(\rbzero.tex_r1[19] ),
    .A2(_04933_),
    .B1(_05212_),
    .C1(_05191_),
    .X(_05213_));
 sky130_fd_sc_hd__a31o_1 _12025_ (.A1(\rbzero.tex_r1[17] ),
    .A2(_04935_),
    .A3(_05186_),
    .B1(_04953_),
    .X(_05214_));
 sky130_fd_sc_hd__a311o_1 _12026_ (.A1(\rbzero.tex_r1[16] ),
    .A2(_04906_),
    .A3(_05181_),
    .B1(_05213_),
    .C1(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__or2_1 _12027_ (.A(\rbzero.tex_r1[30] ),
    .B(_05182_),
    .X(_05216_));
 sky130_fd_sc_hd__o211a_1 _12028_ (.A1(\rbzero.tex_r1[31] ),
    .A2(_05195_),
    .B1(_05216_),
    .C1(_04923_),
    .X(_05217_));
 sky130_fd_sc_hd__a31o_1 _12029_ (.A1(\rbzero.tex_r1[29] ),
    .A2(_05199_),
    .A3(_05032_),
    .B1(_04890_),
    .X(_05218_));
 sky130_fd_sc_hd__a31o_1 _12030_ (.A1(\rbzero.tex_r1[28] ),
    .A2(_05185_),
    .A3(_05195_),
    .B1(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__or2_1 _12031_ (.A(\rbzero.tex_r1[26] ),
    .B(_05032_),
    .X(_05220_));
 sky130_fd_sc_hd__o211a_1 _12032_ (.A1(\rbzero.tex_r1[27] ),
    .A2(_05195_),
    .B1(_05220_),
    .C1(_04923_),
    .X(_05221_));
 sky130_fd_sc_hd__a31o_1 _12033_ (.A1(\rbzero.tex_r1[25] ),
    .A2(_04982_),
    .A3(_05032_),
    .B1(_04919_),
    .X(_05222_));
 sky130_fd_sc_hd__a31o_1 _12034_ (.A1(\rbzero.tex_r1[24] ),
    .A2(_05185_),
    .A3(_05181_),
    .B1(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__o221a_1 _12035_ (.A1(_05217_),
    .A2(_05219_),
    .B1(_05221_),
    .B2(_05223_),
    .C1(_04903_),
    .X(_05224_));
 sky130_fd_sc_hd__a311o_1 _12036_ (.A1(_04955_),
    .A2(_05211_),
    .A3(_05215_),
    .B1(_04887_),
    .C1(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__or2_1 _12037_ (.A(\rbzero.tex_r1[46] ),
    .B(_05031_),
    .X(_05226_));
 sky130_fd_sc_hd__o211a_1 _12038_ (.A1(\rbzero.tex_r1[47] ),
    .A2(_05002_),
    .B1(_05226_),
    .C1(_04922_),
    .X(_05227_));
 sky130_fd_sc_hd__a31o_1 _12039_ (.A1(\rbzero.tex_r1[45] ),
    .A2(_05199_),
    .A3(_05032_),
    .B1(_04890_),
    .X(_05228_));
 sky130_fd_sc_hd__a311o_1 _12040_ (.A1(\rbzero.tex_r1[44] ),
    .A2(_04935_),
    .A3(_05195_),
    .B1(_05227_),
    .C1(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__or2_1 _12041_ (.A(\rbzero.tex_r1[42] ),
    .B(_05031_),
    .X(_05230_));
 sky130_fd_sc_hd__o211a_1 _12042_ (.A1(\rbzero.tex_r1[43] ),
    .A2(_05002_),
    .B1(_05230_),
    .C1(_04922_),
    .X(_05231_));
 sky130_fd_sc_hd__a31o_1 _12043_ (.A1(\rbzero.tex_r1[41] ),
    .A2(_05199_),
    .A3(_05032_),
    .B1(_04952_),
    .X(_05232_));
 sky130_fd_sc_hd__a311o_1 _12044_ (.A1(\rbzero.tex_r1[40] ),
    .A2(_04935_),
    .A3(_05195_),
    .B1(_05231_),
    .C1(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__or2_1 _12045_ (.A(\rbzero.tex_r1[38] ),
    .B(_05031_),
    .X(_05234_));
 sky130_fd_sc_hd__o211a_1 _12046_ (.A1(\rbzero.tex_r1[39] ),
    .A2(_04924_),
    .B1(_05234_),
    .C1(_04944_),
    .X(_05235_));
 sky130_fd_sc_hd__clkbuf_4 _12047_ (.A(_04829_),
    .X(_05236_));
 sky130_fd_sc_hd__a31o_1 _12048_ (.A1(\rbzero.tex_r1[37] ),
    .A2(_05198_),
    .A3(_05236_),
    .B1(_04939_),
    .X(_05237_));
 sky130_fd_sc_hd__a31o_1 _12049_ (.A1(\rbzero.tex_r1[36] ),
    .A2(_04982_),
    .A3(_04924_),
    .B1(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__or2_1 _12050_ (.A(\rbzero.tex_r1[34] ),
    .B(_05236_),
    .X(_05239_));
 sky130_fd_sc_hd__o211a_1 _12051_ (.A1(\rbzero.tex_r1[35] ),
    .A2(_04924_),
    .B1(_05239_),
    .C1(_04944_),
    .X(_05240_));
 sky130_fd_sc_hd__a31o_1 _12052_ (.A1(\rbzero.tex_r1[33] ),
    .A2(_04981_),
    .A3(_05236_),
    .B1(_04918_),
    .X(_05241_));
 sky130_fd_sc_hd__a31o_1 _12053_ (.A1(\rbzero.tex_r1[32] ),
    .A2(_04982_),
    .A3(_04910_),
    .B1(_05241_),
    .X(_05242_));
 sky130_fd_sc_hd__o221a_1 _12054_ (.A1(_05235_),
    .A2(_05238_),
    .B1(_05240_),
    .B2(_05242_),
    .C1(_04967_),
    .X(_05243_));
 sky130_fd_sc_hd__a311o_1 _12055_ (.A1(_04903_),
    .A2(_05229_),
    .A3(_05233_),
    .B1(_04958_),
    .C1(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__or2_1 _12056_ (.A(\rbzero.tex_r1[62] ),
    .B(_05031_),
    .X(_05245_));
 sky130_fd_sc_hd__o211a_1 _12057_ (.A1(\rbzero.tex_r1[63] ),
    .A2(_05002_),
    .B1(_05245_),
    .C1(_04922_),
    .X(_05246_));
 sky130_fd_sc_hd__a31o_1 _12058_ (.A1(\rbzero.tex_r1[61] ),
    .A2(_05199_),
    .A3(_05032_),
    .B1(_04890_),
    .X(_05247_));
 sky130_fd_sc_hd__a311o_1 _12059_ (.A1(\rbzero.tex_r1[60] ),
    .A2(_04935_),
    .A3(_05195_),
    .B1(_05246_),
    .C1(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__or2_1 _12060_ (.A(\rbzero.tex_r1[58] ),
    .B(_05031_),
    .X(_05249_));
 sky130_fd_sc_hd__o211a_1 _12061_ (.A1(\rbzero.tex_r1[59] ),
    .A2(_05002_),
    .B1(_05249_),
    .C1(_04922_),
    .X(_05250_));
 sky130_fd_sc_hd__a31o_1 _12062_ (.A1(\rbzero.tex_r1[57] ),
    .A2(_05199_),
    .A3(_05182_),
    .B1(_04952_),
    .X(_05251_));
 sky130_fd_sc_hd__a311o_1 _12063_ (.A1(\rbzero.tex_r1[56] ),
    .A2(_04935_),
    .A3(_04933_),
    .B1(_05250_),
    .C1(_05251_),
    .X(_05252_));
 sky130_fd_sc_hd__or2_1 _12064_ (.A(\rbzero.tex_r1[54] ),
    .B(_05031_),
    .X(_05253_));
 sky130_fd_sc_hd__o211a_1 _12065_ (.A1(\rbzero.tex_r1[55] ),
    .A2(_04924_),
    .B1(_05253_),
    .C1(_04944_),
    .X(_05254_));
 sky130_fd_sc_hd__a31o_1 _12066_ (.A1(\rbzero.tex_r1[53] ),
    .A2(_05198_),
    .A3(_05236_),
    .B1(_04939_),
    .X(_05255_));
 sky130_fd_sc_hd__a31o_1 _12067_ (.A1(\rbzero.tex_r1[52] ),
    .A2(_05199_),
    .A3(_04924_),
    .B1(_05255_),
    .X(_05256_));
 sky130_fd_sc_hd__or2_1 _12068_ (.A(\rbzero.tex_r1[50] ),
    .B(_05031_),
    .X(_05257_));
 sky130_fd_sc_hd__o211a_1 _12069_ (.A1(\rbzero.tex_r1[51] ),
    .A2(_04924_),
    .B1(_05257_),
    .C1(_04944_),
    .X(_05258_));
 sky130_fd_sc_hd__a31o_1 _12070_ (.A1(\rbzero.tex_r1[49] ),
    .A2(_04981_),
    .A3(_05236_),
    .B1(_04918_),
    .X(_05259_));
 sky130_fd_sc_hd__a31o_1 _12071_ (.A1(\rbzero.tex_r1[48] ),
    .A2(_04982_),
    .A3(_04910_),
    .B1(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__o221a_1 _12072_ (.A1(_05254_),
    .A2(_05256_),
    .B1(_05258_),
    .B2(_05260_),
    .C1(_04967_),
    .X(_05261_));
 sky130_fd_sc_hd__a311o_1 _12073_ (.A1(_04903_),
    .A2(_05248_),
    .A3(_05252_),
    .B1(_04887_),
    .C1(_05261_),
    .X(_05262_));
 sky130_fd_sc_hd__buf_6 _12074_ (.A(net42),
    .X(_05263_));
 sky130_fd_sc_hd__a31o_1 _12075_ (.A1(_04832_),
    .A2(_05244_),
    .A3(_05262_),
    .B1(_05263_),
    .X(_05264_));
 sky130_fd_sc_hd__a31o_1 _12076_ (.A1(_04810_),
    .A2(_05207_),
    .A3(_05225_),
    .B1(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__o211a_1 _12077_ (.A1(_05017_),
    .A2(_05180_),
    .B1(_05265_),
    .C1(_04900_),
    .X(_05266_));
 sky130_fd_sc_hd__mux2_1 _12078_ (.A0(\rbzero.color_sky[1] ),
    .A1(\rbzero.color_floor[1] ),
    .S(_04825_),
    .X(_05267_));
 sky130_fd_sc_hd__and2b_1 _12079_ (.A_N(_04900_),
    .B(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__or4_1 _12080_ (.A(\gpout0.vpos[7] ),
    .B(_04653_),
    .C(_03972_),
    .D(_04410_),
    .X(_05269_));
 sky130_fd_sc_hd__and2_1 _12081_ (.A(_04731_),
    .B(\gpout0.vpos[4] ),
    .X(_05270_));
 sky130_fd_sc_hd__or3b_1 _12082_ (.A(_04672_),
    .B(_04704_),
    .C_N(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__xnor2_1 _12083_ (.A(_04656_),
    .B(_04628_),
    .Y(_05272_));
 sky130_fd_sc_hd__o22ai_1 _12084_ (.A1(_04648_),
    .A2(_04411_),
    .B1(_04578_),
    .B2(_04652_),
    .Y(_05273_));
 sky130_fd_sc_hd__a221o_1 _12085_ (.A1(\gpout0.vpos[4] ),
    .A2(_04418_),
    .B1(_04578_),
    .B2(_04652_),
    .C1(_05273_),
    .X(_05274_));
 sky130_fd_sc_hd__a2bb2o_1 _12086_ (.A1_N(_04651_),
    .A2_N(_04419_),
    .B1(_04411_),
    .B2(_04648_),
    .X(_05275_));
 sky130_fd_sc_hd__or3_1 _12087_ (.A(_05272_),
    .B(_05274_),
    .C(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__o31a_1 _12088_ (.A1(_04579_),
    .A2(_05269_),
    .A3(_05271_),
    .B1(_05276_),
    .X(_05277_));
 sky130_fd_sc_hd__nor2_1 _12089_ (.A(_04741_),
    .B(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__xnor2_1 _12090_ (.A(_04656_),
    .B(_04704_),
    .Y(_05279_));
 sky130_fd_sc_hd__nand2_1 _12091_ (.A(_04654_),
    .B(_04655_),
    .Y(_05280_));
 sky130_fd_sc_hd__nor2_1 _12092_ (.A(_04652_),
    .B(_04412_),
    .Y(_05281_));
 sky130_fd_sc_hd__a31o_1 _12093_ (.A1(_04657_),
    .A2(_04589_),
    .A3(_05280_),
    .B1(_05281_),
    .X(_05282_));
 sky130_fd_sc_hd__and3_1 _12094_ (.A(_03972_),
    .B(_04418_),
    .C(_04411_),
    .X(_05283_));
 sky130_fd_sc_hd__o2bb2a_1 _12095_ (.A1_N(_04415_),
    .A2_N(_05283_),
    .B1(_04700_),
    .B2(_03972_),
    .X(_05284_));
 sky130_fd_sc_hd__a2bb2o_1 _12096_ (.A1_N(\gpout0.vpos[4] ),
    .A2_N(_04578_),
    .B1(_04412_),
    .B2(\gpout0.vpos[3] ),
    .X(_05285_));
 sky130_fd_sc_hd__or4_1 _12097_ (.A(_04648_),
    .B(_04418_),
    .C(_05281_),
    .D(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__a211o_1 _12098_ (.A1(_04651_),
    .A2(_04578_),
    .B1(_05279_),
    .C1(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__or2b_1 _12099_ (.A(_04655_),
    .B_N(_05054_),
    .X(_05288_));
 sky130_fd_sc_hd__o2111a_1 _12100_ (.A1(_04653_),
    .A2(_04695_),
    .B1(_05284_),
    .C1(_05287_),
    .D1(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__a21bo_1 _12101_ (.A1(_05279_),
    .A2(_05282_),
    .B1_N(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__and2_1 _12102_ (.A(_04744_),
    .B(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__o21bai_1 _12103_ (.A1(_04722_),
    .A2(_04729_),
    .B1_N(_04719_),
    .Y(_05292_));
 sky130_fd_sc_hd__a221o_1 _12104_ (.A1(_05278_),
    .A2(_05291_),
    .B1(_05292_),
    .B2(_04744_),
    .C1(_04703_),
    .X(_05293_));
 sky130_fd_sc_hd__o31a_1 _12105_ (.A1(_05047_),
    .A2(_05266_),
    .A3(_05268_),
    .B1(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__nor2_1 _12106_ (.A(_04650_),
    .B(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__o21ai_1 _12107_ (.A1(_05176_),
    .A2(_05295_),
    .B1(_05051_),
    .Y(_05296_));
 sky130_fd_sc_hd__o211ai_4 _12108_ (.A1(_04436_),
    .A2(_04635_),
    .B1(_05056_),
    .C1(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__inv_2 _12109_ (.A(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__mux2_4 _12110_ (.A0(\reg_rgb[7] ),
    .A1(_05298_),
    .S(_05058_),
    .X(_05299_));
 sky130_fd_sc_hd__clkbuf_1 _12111_ (.A(_05299_),
    .X(net69));
 sky130_fd_sc_hd__inv_2 _12112_ (.A(_04650_),
    .Y(_05300_));
 sky130_fd_sc_hd__mux2_1 _12113_ (.A0(\rbzero.tex_g0[7] ),
    .A1(\rbzero.tex_g0[6] ),
    .S(_04933_),
    .X(_05301_));
 sky130_fd_sc_hd__mux2_1 _12114_ (.A0(\rbzero.tex_g0[5] ),
    .A1(\rbzero.tex_g0[4] ),
    .S(_05010_),
    .X(_05302_));
 sky130_fd_sc_hd__or2_1 _12115_ (.A(_05191_),
    .B(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__o211a_1 _12116_ (.A1(_04906_),
    .A2(_05301_),
    .B1(_05303_),
    .C1(_04920_),
    .X(_05304_));
 sky130_fd_sc_hd__buf_4 _12117_ (.A(_05010_),
    .X(_05305_));
 sky130_fd_sc_hd__mux2_1 _12118_ (.A0(\rbzero.tex_g0[1] ),
    .A1(\rbzero.tex_g0[0] ),
    .S(_05305_),
    .X(_05306_));
 sky130_fd_sc_hd__and3_1 _12119_ (.A(\rbzero.tex_g0[3] ),
    .B(_04927_),
    .C(_04929_),
    .X(_05307_));
 sky130_fd_sc_hd__a21o_1 _12120_ (.A1(\rbzero.tex_g0[2] ),
    .A2(_05195_),
    .B1(_05185_),
    .X(_05308_));
 sky130_fd_sc_hd__o221a_1 _12121_ (.A1(_04923_),
    .A2(_05306_),
    .B1(_05307_),
    .B2(_05308_),
    .C1(_04941_),
    .X(_05309_));
 sky130_fd_sc_hd__mux2_1 _12122_ (.A0(\rbzero.tex_g0[9] ),
    .A1(\rbzero.tex_g0[8] ),
    .S(_04932_),
    .X(_05310_));
 sky130_fd_sc_hd__mux2_1 _12123_ (.A0(\rbzero.tex_g0[11] ),
    .A1(\rbzero.tex_g0[10] ),
    .S(_04932_),
    .X(_05311_));
 sky130_fd_sc_hd__mux2_1 _12124_ (.A0(_05310_),
    .A1(_05311_),
    .S(_05191_),
    .X(_05312_));
 sky130_fd_sc_hd__mux2_1 _12125_ (.A0(\rbzero.tex_g0[13] ),
    .A1(\rbzero.tex_g0[12] ),
    .S(_05002_),
    .X(_05313_));
 sky130_fd_sc_hd__buf_4 _12126_ (.A(_04913_),
    .X(_05314_));
 sky130_fd_sc_hd__mux2_1 _12127_ (.A0(\rbzero.tex_g0[15] ),
    .A1(\rbzero.tex_g0[14] ),
    .S(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__or2_1 _12128_ (.A(_04982_),
    .B(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__o211a_1 _12129_ (.A1(_04923_),
    .A2(_05313_),
    .B1(_05316_),
    .C1(_04953_),
    .X(_05317_));
 sky130_fd_sc_hd__a211o_1 _12130_ (.A1(_04941_),
    .A2(_05312_),
    .B1(_05317_),
    .C1(_04955_),
    .X(_05318_));
 sky130_fd_sc_hd__o311a_1 _12131_ (.A1(_04903_),
    .A2(_05304_),
    .A3(_05309_),
    .B1(_05318_),
    .C1(_04887_),
    .X(_05319_));
 sky130_fd_sc_hd__mux2_1 _12132_ (.A0(\rbzero.tex_g0[29] ),
    .A1(\rbzero.tex_g0[28] ),
    .S(_04964_),
    .X(_05320_));
 sky130_fd_sc_hd__mux2_1 _12133_ (.A0(\rbzero.tex_g0[31] ),
    .A1(\rbzero.tex_g0[30] ),
    .S(_05010_),
    .X(_05321_));
 sky130_fd_sc_hd__mux2_1 _12134_ (.A0(_05320_),
    .A1(_05321_),
    .S(_04947_),
    .X(_05322_));
 sky130_fd_sc_hd__mux2_1 _12135_ (.A0(\rbzero.tex_g0[25] ),
    .A1(\rbzero.tex_g0[24] ),
    .S(_05010_),
    .X(_05323_));
 sky130_fd_sc_hd__and3_1 _12136_ (.A(\rbzero.tex_g0[27] ),
    .B(_04927_),
    .C(_04929_),
    .X(_05324_));
 sky130_fd_sc_hd__a21o_1 _12137_ (.A1(\rbzero.tex_g0[26] ),
    .A2(_04924_),
    .B1(_04982_),
    .X(_05325_));
 sky130_fd_sc_hd__o221a_1 _12138_ (.A1(_05191_),
    .A2(_05323_),
    .B1(_05324_),
    .B2(_05325_),
    .C1(_04937_),
    .X(_05326_));
 sky130_fd_sc_hd__a211o_1 _12139_ (.A1(_04920_),
    .A2(_05322_),
    .B1(_05326_),
    .C1(_04955_),
    .X(_05327_));
 sky130_fd_sc_hd__mux2_1 _12140_ (.A0(\rbzero.tex_g0[17] ),
    .A1(\rbzero.tex_g0[16] ),
    .S(_04964_),
    .X(_05328_));
 sky130_fd_sc_hd__mux2_1 _12141_ (.A0(\rbzero.tex_g0[19] ),
    .A1(\rbzero.tex_g0[18] ),
    .S(_05010_),
    .X(_05329_));
 sky130_fd_sc_hd__mux2_1 _12142_ (.A0(_05328_),
    .A1(_05329_),
    .S(_04947_),
    .X(_05330_));
 sky130_fd_sc_hd__mux2_1 _12143_ (.A0(\rbzero.tex_g0[21] ),
    .A1(\rbzero.tex_g0[20] ),
    .S(_04932_),
    .X(_05331_));
 sky130_fd_sc_hd__mux2_1 _12144_ (.A0(\rbzero.tex_g0[23] ),
    .A1(\rbzero.tex_g0[22] ),
    .S(_04931_),
    .X(_05332_));
 sky130_fd_sc_hd__or2_1 _12145_ (.A(_05199_),
    .B(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__o211a_1 _12146_ (.A1(_05191_),
    .A2(_05331_),
    .B1(_05333_),
    .C1(_04953_),
    .X(_05334_));
 sky130_fd_sc_hd__a211o_1 _12147_ (.A1(_04941_),
    .A2(_05330_),
    .B1(_05334_),
    .C1(_04902_),
    .X(_05335_));
 sky130_fd_sc_hd__a31o_1 _12148_ (.A1(_04958_),
    .A2(_05327_),
    .A3(_05335_),
    .B1(_04832_),
    .X(_05336_));
 sky130_fd_sc_hd__mux2_1 _12149_ (.A0(\rbzero.tex_g0[39] ),
    .A1(\rbzero.tex_g0[38] ),
    .S(_05010_),
    .X(_05337_));
 sky130_fd_sc_hd__mux2_1 _12150_ (.A0(\rbzero.tex_g0[37] ),
    .A1(\rbzero.tex_g0[36] ),
    .S(_04948_),
    .X(_05338_));
 sky130_fd_sc_hd__mux2_1 _12151_ (.A0(_05337_),
    .A1(_05338_),
    .S(_04935_),
    .X(_05339_));
 sky130_fd_sc_hd__mux2_1 _12152_ (.A0(\rbzero.tex_g0[33] ),
    .A1(\rbzero.tex_g0[32] ),
    .S(_05010_),
    .X(_05340_));
 sky130_fd_sc_hd__mux2_1 _12153_ (.A0(\rbzero.tex_g0[35] ),
    .A1(\rbzero.tex_g0[34] ),
    .S(_04948_),
    .X(_05341_));
 sky130_fd_sc_hd__mux2_1 _12154_ (.A0(_05340_),
    .A1(_05341_),
    .S(_04912_),
    .X(_05342_));
 sky130_fd_sc_hd__mux2_1 _12155_ (.A0(_05339_),
    .A1(_05342_),
    .S(_04941_),
    .X(_05343_));
 sky130_fd_sc_hd__mux2_1 _12156_ (.A0(\rbzero.tex_g0[47] ),
    .A1(\rbzero.tex_g0[46] ),
    .S(_04933_),
    .X(_05344_));
 sky130_fd_sc_hd__mux2_1 _12157_ (.A0(\rbzero.tex_g0[45] ),
    .A1(\rbzero.tex_g0[44] ),
    .S(_05002_),
    .X(_05345_));
 sky130_fd_sc_hd__or2_1 _12158_ (.A(_04923_),
    .B(_05345_),
    .X(_05346_));
 sky130_fd_sc_hd__o211a_1 _12159_ (.A1(_04906_),
    .A2(_05344_),
    .B1(_05346_),
    .C1(_04920_),
    .X(_05347_));
 sky130_fd_sc_hd__mux2_1 _12160_ (.A0(\rbzero.tex_g0[41] ),
    .A1(\rbzero.tex_g0[40] ),
    .S(_05002_),
    .X(_05348_));
 sky130_fd_sc_hd__mux2_1 _12161_ (.A0(\rbzero.tex_g0[43] ),
    .A1(\rbzero.tex_g0[42] ),
    .S(_04932_),
    .X(_05349_));
 sky130_fd_sc_hd__mux2_1 _12162_ (.A0(_05348_),
    .A1(_05349_),
    .S(_05191_),
    .X(_05350_));
 sky130_fd_sc_hd__a21o_1 _12163_ (.A1(_04941_),
    .A2(_05350_),
    .B1(_04955_),
    .X(_05351_));
 sky130_fd_sc_hd__o221a_1 _12164_ (.A1(_04903_),
    .A2(_05343_),
    .B1(_05347_),
    .B2(_05351_),
    .C1(_04887_),
    .X(_05352_));
 sky130_fd_sc_hd__mux2_1 _12165_ (.A0(\rbzero.tex_g0[53] ),
    .A1(\rbzero.tex_g0[52] ),
    .S(_04932_),
    .X(_05353_));
 sky130_fd_sc_hd__mux2_1 _12166_ (.A0(\rbzero.tex_g0[55] ),
    .A1(\rbzero.tex_g0[54] ),
    .S(_04964_),
    .X(_05354_));
 sky130_fd_sc_hd__mux2_1 _12167_ (.A0(_05353_),
    .A1(_05354_),
    .S(_05191_),
    .X(_05355_));
 sky130_fd_sc_hd__mux2_1 _12168_ (.A0(\rbzero.tex_g0[49] ),
    .A1(\rbzero.tex_g0[48] ),
    .S(_04964_),
    .X(_05356_));
 sky130_fd_sc_hd__and3_1 _12169_ (.A(\rbzero.tex_g0[51] ),
    .B(_04927_),
    .C(_04929_),
    .X(_05357_));
 sky130_fd_sc_hd__a21o_1 _12170_ (.A1(\rbzero.tex_g0[50] ),
    .A2(_04924_),
    .B1(_04982_),
    .X(_05358_));
 sky130_fd_sc_hd__o221a_1 _12171_ (.A1(_05191_),
    .A2(_05356_),
    .B1(_05357_),
    .B2(_05358_),
    .C1(_04937_),
    .X(_05359_));
 sky130_fd_sc_hd__a211o_1 _12172_ (.A1(_04920_),
    .A2(_05355_),
    .B1(_05359_),
    .C1(_04903_),
    .X(_05360_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(\rbzero.tex_g0[57] ),
    .A1(\rbzero.tex_g0[56] ),
    .S(_04932_),
    .X(_05361_));
 sky130_fd_sc_hd__mux2_1 _12174_ (.A0(\rbzero.tex_g0[59] ),
    .A1(\rbzero.tex_g0[58] ),
    .S(_04964_),
    .X(_05362_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(_05361_),
    .A1(_05362_),
    .S(_04947_),
    .X(_05363_));
 sky130_fd_sc_hd__and2_1 _12176_ (.A(\rbzero.tex_g0[62] ),
    .B(_05002_),
    .X(_05364_));
 sky130_fd_sc_hd__a31o_1 _12177_ (.A1(\rbzero.tex_g0[63] ),
    .A2(_04927_),
    .A3(_04929_),
    .B1(_05199_),
    .X(_05365_));
 sky130_fd_sc_hd__mux2_1 _12178_ (.A0(\rbzero.tex_g0[61] ),
    .A1(\rbzero.tex_g0[60] ),
    .S(_04932_),
    .X(_05366_));
 sky130_fd_sc_hd__o221a_1 _12179_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05366_),
    .B2(_05191_),
    .C1(_04953_),
    .X(_05367_));
 sky130_fd_sc_hd__a211o_1 _12180_ (.A1(_04941_),
    .A2(_05363_),
    .B1(_05367_),
    .C1(_04955_),
    .X(_05368_));
 sky130_fd_sc_hd__a31o_1 _12181_ (.A1(_04958_),
    .A2(_05360_),
    .A3(_05368_),
    .B1(_04810_),
    .X(_05369_));
 sky130_fd_sc_hd__o221a_2 _12182_ (.A1(_05319_),
    .A2(_05336_),
    .B1(_05352_),
    .B2(_05369_),
    .C1(_05017_),
    .X(_05370_));
 sky130_fd_sc_hd__or3b_1 _12183_ (.A(_05027_),
    .B(_05026_),
    .C_N(\rbzero.row_render.wall[0] ),
    .X(_05371_));
 sky130_fd_sc_hd__or3_1 _12184_ (.A(_04890_),
    .B(_04934_),
    .C(_05002_),
    .X(_05372_));
 sky130_fd_sc_hd__or2b_1 _12185_ (.A(_05372_),
    .B_N(_05036_),
    .X(_05373_));
 sky130_fd_sc_hd__a311o_1 _12186_ (.A1(\rbzero.row_render.side ),
    .A2(_05033_),
    .A3(_05373_),
    .B1(_05038_),
    .C1(_05020_),
    .X(_05374_));
 sky130_fd_sc_hd__a31o_1 _12187_ (.A1(_05019_),
    .A2(_05371_),
    .A3(_05374_),
    .B1(_05043_),
    .X(_05375_));
 sky130_fd_sc_hd__nand2_1 _12188_ (.A(_04900_),
    .B(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__mux2_1 _12189_ (.A0(\rbzero.color_sky[2] ),
    .A1(\rbzero.color_floor[2] ),
    .S(_04825_),
    .X(_05377_));
 sky130_fd_sc_hd__o221ai_2 _12190_ (.A1(_05370_),
    .A2(_05376_),
    .B1(_05377_),
    .B2(_04900_),
    .C1(_04702_),
    .Y(_05378_));
 sky130_fd_sc_hd__nand2_1 _12191_ (.A(_05047_),
    .B(_04683_),
    .Y(_05379_));
 sky130_fd_sc_hd__a31o_1 _12192_ (.A1(_05300_),
    .A2(_05378_),
    .A3(_05379_),
    .B1(_04661_),
    .X(_05380_));
 sky130_fd_sc_hd__nand2_1 _12193_ (.A(_05051_),
    .B(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__o211a_4 _12194_ (.A1(_04429_),
    .A2(_04635_),
    .B1(_05056_),
    .C1(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__mux2_2 _12195_ (.A0(\reg_rgb[14] ),
    .A1(_05382_),
    .S(_05058_),
    .X(_05383_));
 sky130_fd_sc_hd__clkbuf_1 _12196_ (.A(_05383_),
    .X(net64));
 sky130_fd_sc_hd__or2_1 _12197_ (.A(\rbzero.tex_g1[14] ),
    .B(_05236_),
    .X(_05384_));
 sky130_fd_sc_hd__o211a_1 _12198_ (.A1(\rbzero.tex_g1[15] ),
    .A2(_04910_),
    .B1(_05384_),
    .C1(_04912_),
    .X(_05385_));
 sky130_fd_sc_hd__a31o_1 _12199_ (.A1(\rbzero.tex_g1[13] ),
    .A2(_04905_),
    .A3(_05186_),
    .B1(_04940_),
    .X(_05386_));
 sky130_fd_sc_hd__a311o_1 _12200_ (.A1(\rbzero.tex_g1[12] ),
    .A2(_04906_),
    .A3(_05181_),
    .B1(_05385_),
    .C1(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__or2_1 _12201_ (.A(\rbzero.tex_g1[10] ),
    .B(_05236_),
    .X(_05388_));
 sky130_fd_sc_hd__o211a_1 _12202_ (.A1(\rbzero.tex_g1[11] ),
    .A2(_04910_),
    .B1(_05388_),
    .C1(_04912_),
    .X(_05389_));
 sky130_fd_sc_hd__a31o_1 _12203_ (.A1(\rbzero.tex_g1[9] ),
    .A2(_04905_),
    .A3(_05186_),
    .B1(_04919_),
    .X(_05390_));
 sky130_fd_sc_hd__a311o_1 _12204_ (.A1(\rbzero.tex_g1[8] ),
    .A2(_04906_),
    .A3(_05181_),
    .B1(_05389_),
    .C1(_05390_),
    .X(_05391_));
 sky130_fd_sc_hd__or2_1 _12205_ (.A(\rbzero.tex_g1[6] ),
    .B(_04831_),
    .X(_05392_));
 sky130_fd_sc_hd__o211a_1 _12206_ (.A1(\rbzero.tex_g1[7] ),
    .A2(_05305_),
    .B1(_05392_),
    .C1(_04947_),
    .X(_05393_));
 sky130_fd_sc_hd__a31o_1 _12207_ (.A1(\rbzero.tex_g1[5] ),
    .A2(_04981_),
    .A3(_04831_),
    .B1(_04939_),
    .X(_05394_));
 sky130_fd_sc_hd__a31o_1 _12208_ (.A1(\rbzero.tex_g1[4] ),
    .A2(_04935_),
    .A3(_05305_),
    .B1(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__or2_1 _12209_ (.A(\rbzero.tex_g1[2] ),
    .B(_04831_),
    .X(_05396_));
 sky130_fd_sc_hd__o211a_1 _12210_ (.A1(\rbzero.tex_g1[3] ),
    .A2(_05305_),
    .B1(_05396_),
    .C1(_04947_),
    .X(_05397_));
 sky130_fd_sc_hd__a31o_1 _12211_ (.A1(\rbzero.tex_g1[1] ),
    .A2(_04904_),
    .A3(_05182_),
    .B1(_04918_),
    .X(_05398_));
 sky130_fd_sc_hd__a31o_1 _12212_ (.A1(\rbzero.tex_g1[0] ),
    .A2(_04935_),
    .A3(_04933_),
    .B1(_05398_),
    .X(_05399_));
 sky130_fd_sc_hd__o221a_1 _12213_ (.A1(_05393_),
    .A2(_05395_),
    .B1(_05397_),
    .B2(_05399_),
    .C1(_04967_),
    .X(_05400_));
 sky130_fd_sc_hd__a311o_1 _12214_ (.A1(_04903_),
    .A2(_05387_),
    .A3(_05391_),
    .B1(_04958_),
    .C1(_05400_),
    .X(_05401_));
 sky130_fd_sc_hd__or2_1 _12215_ (.A(\rbzero.tex_g1[22] ),
    .B(_05236_),
    .X(_05402_));
 sky130_fd_sc_hd__o211a_1 _12216_ (.A1(\rbzero.tex_g1[23] ),
    .A2(_04910_),
    .B1(_05402_),
    .C1(_04912_),
    .X(_05403_));
 sky130_fd_sc_hd__a31o_1 _12217_ (.A1(\rbzero.tex_g1[21] ),
    .A2(_04905_),
    .A3(_05186_),
    .B1(_04940_),
    .X(_05404_));
 sky130_fd_sc_hd__a311o_1 _12218_ (.A1(\rbzero.tex_g1[20] ),
    .A2(_05185_),
    .A3(_05181_),
    .B1(_05403_),
    .C1(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__or2_1 _12219_ (.A(\rbzero.tex_g1[18] ),
    .B(_05236_),
    .X(_05406_));
 sky130_fd_sc_hd__o211a_1 _12220_ (.A1(\rbzero.tex_g1[19] ),
    .A2(_04910_),
    .B1(_05406_),
    .C1(_04912_),
    .X(_05407_));
 sky130_fd_sc_hd__a31o_1 _12221_ (.A1(\rbzero.tex_g1[17] ),
    .A2(_04905_),
    .A3(_05186_),
    .B1(_04919_),
    .X(_05408_));
 sky130_fd_sc_hd__a311o_1 _12222_ (.A1(\rbzero.tex_g1[16] ),
    .A2(_05185_),
    .A3(_05181_),
    .B1(_05407_),
    .C1(_05408_),
    .X(_05409_));
 sky130_fd_sc_hd__or2_1 _12223_ (.A(\rbzero.tex_g1[30] ),
    .B(_05236_),
    .X(_05410_));
 sky130_fd_sc_hd__o211a_1 _12224_ (.A1(\rbzero.tex_g1[31] ),
    .A2(_05305_),
    .B1(_05410_),
    .C1(_04912_),
    .X(_05411_));
 sky130_fd_sc_hd__a31o_1 _12225_ (.A1(\rbzero.tex_g1[29] ),
    .A2(_04981_),
    .A3(_04831_),
    .B1(_04939_),
    .X(_05412_));
 sky130_fd_sc_hd__a31o_1 _12226_ (.A1(\rbzero.tex_g1[28] ),
    .A2(_04905_),
    .A3(_05305_),
    .B1(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__or2_1 _12227_ (.A(\rbzero.tex_g1[26] ),
    .B(_04831_),
    .X(_05414_));
 sky130_fd_sc_hd__o211a_1 _12228_ (.A1(\rbzero.tex_g1[27] ),
    .A2(_05305_),
    .B1(_05414_),
    .C1(_04947_),
    .X(_05415_));
 sky130_fd_sc_hd__a31o_1 _12229_ (.A1(\rbzero.tex_g1[25] ),
    .A2(_04904_),
    .A3(_05182_),
    .B1(_04918_),
    .X(_05416_));
 sky130_fd_sc_hd__a31o_1 _12230_ (.A1(\rbzero.tex_g1[24] ),
    .A2(_04935_),
    .A3(_04933_),
    .B1(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__o221a_1 _12231_ (.A1(_05411_),
    .A2(_05413_),
    .B1(_05415_),
    .B2(_05417_),
    .C1(_04902_),
    .X(_05418_));
 sky130_fd_sc_hd__a311o_1 _12232_ (.A1(_04955_),
    .A2(_05405_),
    .A3(_05409_),
    .B1(_04887_),
    .C1(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__or2_1 _12233_ (.A(\rbzero.tex_g1[54] ),
    .B(_04830_),
    .X(_05420_));
 sky130_fd_sc_hd__o211a_1 _12234_ (.A1(\rbzero.tex_g1[55] ),
    .A2(_04948_),
    .B1(_05420_),
    .C1(_04827_),
    .X(_05421_));
 sky130_fd_sc_hd__a31o_1 _12235_ (.A1(\rbzero.tex_g1[53] ),
    .A2(_04904_),
    .A3(_05182_),
    .B1(_04939_),
    .X(_05422_));
 sky130_fd_sc_hd__a311o_1 _12236_ (.A1(\rbzero.tex_g1[52] ),
    .A2(_04905_),
    .A3(_05305_),
    .B1(_05421_),
    .C1(_05422_),
    .X(_05423_));
 sky130_fd_sc_hd__or2_1 _12237_ (.A(\rbzero.tex_g1[50] ),
    .B(_04829_),
    .X(_05424_));
 sky130_fd_sc_hd__o211a_1 _12238_ (.A1(\rbzero.tex_g1[51] ),
    .A2(_04948_),
    .B1(_05424_),
    .C1(_04827_),
    .X(_05425_));
 sky130_fd_sc_hd__a31o_1 _12239_ (.A1(\rbzero.tex_g1[49] ),
    .A2(_04904_),
    .A3(_04831_),
    .B1(_04918_),
    .X(_05426_));
 sky130_fd_sc_hd__a311o_1 _12240_ (.A1(\rbzero.tex_g1[48] ),
    .A2(_04905_),
    .A3(_05305_),
    .B1(_05425_),
    .C1(_05426_),
    .X(_05427_));
 sky130_fd_sc_hd__or2_1 _12241_ (.A(\rbzero.tex_g1[62] ),
    .B(_04830_),
    .X(_05428_));
 sky130_fd_sc_hd__o211a_1 _12242_ (.A1(\rbzero.tex_g1[63] ),
    .A2(_05010_),
    .B1(_05428_),
    .C1(_04946_),
    .X(_05429_));
 sky130_fd_sc_hd__a31o_1 _12243_ (.A1(\rbzero.tex_g1[61] ),
    .A2(_04891_),
    .A3(_04830_),
    .B1(_04814_),
    .X(_05430_));
 sky130_fd_sc_hd__a31o_1 _12244_ (.A1(\rbzero.tex_g1[60] ),
    .A2(_04904_),
    .A3(_04964_),
    .B1(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__or2_1 _12245_ (.A(\rbzero.tex_g1[58] ),
    .B(_04830_),
    .X(_05432_));
 sky130_fd_sc_hd__o211a_1 _12246_ (.A1(\rbzero.tex_g1[59] ),
    .A2(_04964_),
    .B1(_05432_),
    .C1(_04946_),
    .X(_05433_));
 sky130_fd_sc_hd__a31o_1 _12247_ (.A1(\rbzero.tex_g1[57] ),
    .A2(_04891_),
    .A3(_05031_),
    .B1(_04917_),
    .X(_05434_));
 sky130_fd_sc_hd__a31o_1 _12248_ (.A1(\rbzero.tex_g1[56] ),
    .A2(_04934_),
    .A3(_04932_),
    .B1(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__o221a_1 _12249_ (.A1(_05429_),
    .A2(_05431_),
    .B1(_05433_),
    .B2(_05435_),
    .C1(_04812_),
    .X(_05436_));
 sky130_fd_sc_hd__a311o_1 _12250_ (.A1(_04967_),
    .A2(_05423_),
    .A3(_05427_),
    .B1(_04887_),
    .C1(_05436_),
    .X(_05437_));
 sky130_fd_sc_hd__or2_1 _12251_ (.A(\rbzero.tex_g1[46] ),
    .B(_04829_),
    .X(_05438_));
 sky130_fd_sc_hd__o211a_1 _12252_ (.A1(\rbzero.tex_g1[47] ),
    .A2(_04948_),
    .B1(_05438_),
    .C1(_04827_),
    .X(_05439_));
 sky130_fd_sc_hd__a31o_1 _12253_ (.A1(\rbzero.tex_g1[45] ),
    .A2(_04904_),
    .A3(_04831_),
    .B1(_04939_),
    .X(_05440_));
 sky130_fd_sc_hd__a311o_1 _12254_ (.A1(\rbzero.tex_g1[44] ),
    .A2(_04905_),
    .A3(_05305_),
    .B1(_05439_),
    .C1(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__or2_1 _12255_ (.A(\rbzero.tex_g1[42] ),
    .B(_04829_),
    .X(_05442_));
 sky130_fd_sc_hd__o211a_1 _12256_ (.A1(\rbzero.tex_g1[43] ),
    .A2(_04948_),
    .B1(_05442_),
    .C1(_04827_),
    .X(_05443_));
 sky130_fd_sc_hd__a31o_1 _12257_ (.A1(\rbzero.tex_g1[41] ),
    .A2(_04904_),
    .A3(_04831_),
    .B1(_04918_),
    .X(_05444_));
 sky130_fd_sc_hd__a311o_1 _12258_ (.A1(\rbzero.tex_g1[40] ),
    .A2(_04905_),
    .A3(_04910_),
    .B1(_05443_),
    .C1(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__or2_1 _12259_ (.A(\rbzero.tex_g1[38] ),
    .B(_04830_),
    .X(_05446_));
 sky130_fd_sc_hd__o211a_1 _12260_ (.A1(\rbzero.tex_g1[39] ),
    .A2(_05010_),
    .B1(_05446_),
    .C1(_04946_),
    .X(_05447_));
 sky130_fd_sc_hd__a31o_1 _12261_ (.A1(\rbzero.tex_g1[37] ),
    .A2(_04817_),
    .A3(_04830_),
    .B1(_04814_),
    .X(_05448_));
 sky130_fd_sc_hd__a31o_1 _12262_ (.A1(\rbzero.tex_g1[36] ),
    .A2(_04904_),
    .A3(_04964_),
    .B1(_05448_),
    .X(_05449_));
 sky130_fd_sc_hd__or2_1 _12263_ (.A(\rbzero.tex_g1[34] ),
    .B(_04830_),
    .X(_05450_));
 sky130_fd_sc_hd__o211a_1 _12264_ (.A1(\rbzero.tex_g1[35] ),
    .A2(_04964_),
    .B1(_05450_),
    .C1(_04946_),
    .X(_05451_));
 sky130_fd_sc_hd__a31o_1 _12265_ (.A1(\rbzero.tex_g1[33] ),
    .A2(_04891_),
    .A3(_04830_),
    .B1(_04917_),
    .X(_05452_));
 sky130_fd_sc_hd__a31o_1 _12266_ (.A1(\rbzero.tex_g1[32] ),
    .A2(_04934_),
    .A3(_04932_),
    .B1(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__o221a_1 _12267_ (.A1(_05447_),
    .A2(_05449_),
    .B1(_05451_),
    .B2(_05453_),
    .C1(_04889_),
    .X(_05454_));
 sky130_fd_sc_hd__a311o_1 _12268_ (.A1(_04902_),
    .A2(_05441_),
    .A3(_05445_),
    .B1(_04823_),
    .C1(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__a31o_1 _12269_ (.A1(_04832_),
    .A2(_05437_),
    .A3(_05455_),
    .B1(net42),
    .X(_05456_));
 sky130_fd_sc_hd__a31oi_4 _12270_ (.A1(_04810_),
    .A2(_05401_),
    .A3(_05419_),
    .B1(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__nand2_1 _12271_ (.A(\rbzero.row_render.side ),
    .B(_05037_),
    .Y(_05458_));
 sky130_fd_sc_hd__a21oi_1 _12272_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_04920_),
    .B1(_05019_),
    .Y(_05459_));
 sky130_fd_sc_hd__o21ai_1 _12273_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_04920_),
    .B1(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__o211a_1 _12274_ (.A1(_05020_),
    .A2(_05458_),
    .B1(_05460_),
    .C1(_05263_),
    .X(_05461_));
 sky130_fd_sc_hd__or3b_1 _12275_ (.A(_05457_),
    .B(_05461_),
    .C_N(_04900_),
    .X(_05462_));
 sky130_fd_sc_hd__mux2_1 _12276_ (.A0(\rbzero.color_sky[3] ),
    .A1(\rbzero.color_floor[3] ),
    .S(_04825_),
    .X(_05463_));
 sky130_fd_sc_hd__or2b_1 _12277_ (.A(_04900_),
    .B_N(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__nor2_1 _12278_ (.A(_04741_),
    .B(_05292_),
    .Y(_05465_));
 sky130_fd_sc_hd__a31oi_1 _12279_ (.A1(_05277_),
    .A2(_05291_),
    .A3(_05465_),
    .B1(_04703_),
    .Y(_05466_));
 sky130_fd_sc_hd__a31oi_1 _12280_ (.A1(_04702_),
    .A2(_05462_),
    .A3(_05464_),
    .B1(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__nor2_1 _12281_ (.A(_04650_),
    .B(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__o21ai_1 _12282_ (.A1(_05176_),
    .A2(_05468_),
    .B1(_05051_),
    .Y(_05469_));
 sky130_fd_sc_hd__o211a_2 _12283_ (.A1(\rbzero.trace_state[3] ),
    .A2(_04635_),
    .B1(_05056_),
    .C1(_05469_),
    .X(_05470_));
 sky130_fd_sc_hd__mux2_2 _12284_ (.A0(\reg_rgb[15] ),
    .A1(_05470_),
    .S(_05058_),
    .X(_05471_));
 sky130_fd_sc_hd__clkbuf_1 _12285_ (.A(_05471_),
    .X(net65));
 sky130_fd_sc_hd__mux2_1 _12286_ (.A0(\rbzero.color_sky[4] ),
    .A1(\rbzero.color_floor[4] ),
    .S(_04825_),
    .X(_05472_));
 sky130_fd_sc_hd__mux2_1 _12287_ (.A0(\rbzero.tex_b0[57] ),
    .A1(\rbzero.tex_b0[56] ),
    .S(_05009_),
    .X(_05473_));
 sky130_fd_sc_hd__mux2_1 _12288_ (.A0(\rbzero.tex_b0[59] ),
    .A1(\rbzero.tex_b0[58] ),
    .S(_05009_),
    .X(_05474_));
 sky130_fd_sc_hd__mux2_1 _12289_ (.A0(_05473_),
    .A1(_05474_),
    .S(_04946_),
    .X(_05475_));
 sky130_fd_sc_hd__and3_1 _12290_ (.A(\rbzero.tex_b0[63] ),
    .B(_04926_),
    .C(_04928_),
    .X(_05476_));
 sky130_fd_sc_hd__a21o_1 _12291_ (.A1(\rbzero.tex_b0[62] ),
    .A2(_04978_),
    .B1(_05198_),
    .X(_05477_));
 sky130_fd_sc_hd__mux2_1 _12292_ (.A0(\rbzero.tex_b0[61] ),
    .A1(\rbzero.tex_b0[60] ),
    .S(_05009_),
    .X(_05478_));
 sky130_fd_sc_hd__o221a_1 _12293_ (.A1(_05476_),
    .A2(_05477_),
    .B1(_05478_),
    .B2(_05190_),
    .C1(_04952_),
    .X(_05479_));
 sky130_fd_sc_hd__a211o_1 _12294_ (.A1(_04937_),
    .A2(_05475_),
    .B1(_05479_),
    .C1(_04967_),
    .X(_05480_));
 sky130_fd_sc_hd__mux2_1 _12295_ (.A0(\rbzero.tex_b0[49] ),
    .A1(\rbzero.tex_b0[48] ),
    .S(_05009_),
    .X(_05481_));
 sky130_fd_sc_hd__mux2_1 _12296_ (.A0(\rbzero.tex_b0[51] ),
    .A1(\rbzero.tex_b0[50] ),
    .S(_04908_),
    .X(_05482_));
 sky130_fd_sc_hd__mux2_1 _12297_ (.A0(_05481_),
    .A1(_05482_),
    .S(_04946_),
    .X(_05483_));
 sky130_fd_sc_hd__and2_1 _12298_ (.A(\rbzero.tex_b0[54] ),
    .B(_05314_),
    .X(_05484_));
 sky130_fd_sc_hd__a31o_1 _12299_ (.A1(\rbzero.tex_b0[55] ),
    .A2(_04926_),
    .A3(_04928_),
    .B1(_04891_),
    .X(_05485_));
 sky130_fd_sc_hd__mux2_1 _12300_ (.A0(\rbzero.tex_b0[53] ),
    .A1(\rbzero.tex_b0[52] ),
    .S(_05009_),
    .X(_05486_));
 sky130_fd_sc_hd__o221a_1 _12301_ (.A1(_05484_),
    .A2(_05485_),
    .B1(_05486_),
    .B2(_05190_),
    .C1(_04952_),
    .X(_05487_));
 sky130_fd_sc_hd__a211o_1 _12302_ (.A1(_04937_),
    .A2(_05483_),
    .B1(_05487_),
    .C1(_04902_),
    .X(_05488_));
 sky130_fd_sc_hd__and3_1 _12303_ (.A(\rbzero.tex_b0[35] ),
    .B(_04926_),
    .C(_04928_),
    .X(_05489_));
 sky130_fd_sc_hd__a21o_1 _12304_ (.A1(\rbzero.tex_b0[34] ),
    .A2(_05314_),
    .B1(_04891_),
    .X(_05490_));
 sky130_fd_sc_hd__mux2_1 _12305_ (.A0(\rbzero.tex_b0[33] ),
    .A1(\rbzero.tex_b0[32] ),
    .S(_04908_),
    .X(_05491_));
 sky130_fd_sc_hd__o221a_1 _12306_ (.A1(_05489_),
    .A2(_05490_),
    .B1(_05491_),
    .B2(_04946_),
    .C1(_04890_),
    .X(_05492_));
 sky130_fd_sc_hd__mux2_1 _12307_ (.A0(\rbzero.tex_b0[37] ),
    .A1(\rbzero.tex_b0[36] ),
    .S(_04908_),
    .X(_05493_));
 sky130_fd_sc_hd__and2_1 _12308_ (.A(\rbzero.tex_b0[38] ),
    .B(_05314_),
    .X(_05494_));
 sky130_fd_sc_hd__a31o_1 _12309_ (.A1(\rbzero.tex_b0[39] ),
    .A2(_04926_),
    .A3(_04928_),
    .B1(_05198_),
    .X(_05495_));
 sky130_fd_sc_hd__o221a_1 _12310_ (.A1(_04946_),
    .A2(_05493_),
    .B1(_05494_),
    .B2(_05495_),
    .C1(_04952_),
    .X(_05496_));
 sky130_fd_sc_hd__mux2_1 _12311_ (.A0(\rbzero.tex_b0[47] ),
    .A1(\rbzero.tex_b0[46] ),
    .S(_04893_),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _12312_ (.A0(\rbzero.tex_b0[45] ),
    .A1(\rbzero.tex_b0[44] ),
    .S(_04907_),
    .X(_05498_));
 sky130_fd_sc_hd__mux2_1 _12313_ (.A0(_05497_),
    .A1(_05498_),
    .S(_04891_),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_1 _12314_ (.A0(\rbzero.tex_b0[41] ),
    .A1(\rbzero.tex_b0[40] ),
    .S(_04907_),
    .X(_05500_));
 sky130_fd_sc_hd__and3_1 _12315_ (.A(\rbzero.tex_b0[43] ),
    .B(_04926_),
    .C(_04928_),
    .X(_05501_));
 sky130_fd_sc_hd__a21o_1 _12316_ (.A1(\rbzero.tex_b0[42] ),
    .A2(_04913_),
    .B1(_04817_),
    .X(_05502_));
 sky130_fd_sc_hd__o221a_1 _12317_ (.A1(_04826_),
    .A2(_05500_),
    .B1(_05501_),
    .B2(_05502_),
    .C1(_04939_),
    .X(_05503_));
 sky130_fd_sc_hd__a211o_1 _12318_ (.A1(_04952_),
    .A2(_05499_),
    .B1(_05503_),
    .C1(_04889_),
    .X(_05504_));
 sky130_fd_sc_hd__o311a_1 _12319_ (.A1(_04812_),
    .A2(_05492_),
    .A3(_05496_),
    .B1(_05504_),
    .C1(_04886_),
    .X(_05505_));
 sky130_fd_sc_hd__a311o_1 _12320_ (.A1(_04958_),
    .A2(_05480_),
    .A3(_05488_),
    .B1(_05505_),
    .C1(_04810_),
    .X(_05506_));
 sky130_fd_sc_hd__mux2_1 _12321_ (.A0(\rbzero.tex_b0[31] ),
    .A1(\rbzero.tex_b0[30] ),
    .S(_05009_),
    .X(_05507_));
 sky130_fd_sc_hd__mux2_1 _12322_ (.A0(\rbzero.tex_b0[29] ),
    .A1(\rbzero.tex_b0[28] ),
    .S(_05009_),
    .X(_05508_));
 sky130_fd_sc_hd__mux2_1 _12323_ (.A0(_05507_),
    .A1(_05508_),
    .S(_04934_),
    .X(_05509_));
 sky130_fd_sc_hd__mux2_1 _12324_ (.A0(\rbzero.tex_b0[25] ),
    .A1(\rbzero.tex_b0[24] ),
    .S(_04908_),
    .X(_05510_));
 sky130_fd_sc_hd__and2_1 _12325_ (.A(\rbzero.tex_b0[26] ),
    .B(_04978_),
    .X(_05511_));
 sky130_fd_sc_hd__a31o_1 _12326_ (.A1(\rbzero.tex_b0[27] ),
    .A2(_04926_),
    .A3(_04928_),
    .B1(_05198_),
    .X(_05512_));
 sky130_fd_sc_hd__o221a_1 _12327_ (.A1(_05190_),
    .A2(_05510_),
    .B1(_05511_),
    .B2(_05512_),
    .C1(_04890_),
    .X(_05513_));
 sky130_fd_sc_hd__a211o_1 _12328_ (.A1(_04953_),
    .A2(_05509_),
    .B1(_05513_),
    .C1(_04967_),
    .X(_05514_));
 sky130_fd_sc_hd__mux2_1 _12329_ (.A0(\rbzero.tex_b0[23] ),
    .A1(\rbzero.tex_b0[22] ),
    .S(_05009_),
    .X(_05515_));
 sky130_fd_sc_hd__mux2_1 _12330_ (.A0(\rbzero.tex_b0[21] ),
    .A1(\rbzero.tex_b0[20] ),
    .S(_04908_),
    .X(_05516_));
 sky130_fd_sc_hd__mux2_1 _12331_ (.A0(_05515_),
    .A1(_05516_),
    .S(_04934_),
    .X(_05517_));
 sky130_fd_sc_hd__mux2_1 _12332_ (.A0(\rbzero.tex_b0[17] ),
    .A1(\rbzero.tex_b0[16] ),
    .S(_04908_),
    .X(_05518_));
 sky130_fd_sc_hd__and2_1 _12333_ (.A(\rbzero.tex_b0[18] ),
    .B(_05314_),
    .X(_05519_));
 sky130_fd_sc_hd__a31o_1 _12334_ (.A1(\rbzero.tex_b0[19] ),
    .A2(_04926_),
    .A3(_04928_),
    .B1(_05198_),
    .X(_05520_));
 sky130_fd_sc_hd__o221a_1 _12335_ (.A1(_04946_),
    .A2(_05518_),
    .B1(_05519_),
    .B2(_05520_),
    .C1(_04890_),
    .X(_05521_));
 sky130_fd_sc_hd__a211o_1 _12336_ (.A1(_04953_),
    .A2(_05517_),
    .B1(_05521_),
    .C1(_04812_),
    .X(_05522_));
 sky130_fd_sc_hd__mux2_1 _12337_ (.A0(\rbzero.tex_b0[3] ),
    .A1(\rbzero.tex_b0[2] ),
    .S(_04907_),
    .X(_05523_));
 sky130_fd_sc_hd__mux2_1 _12338_ (.A0(\rbzero.tex_b0[1] ),
    .A1(\rbzero.tex_b0[0] ),
    .S(_04907_),
    .X(_05524_));
 sky130_fd_sc_hd__mux2_1 _12339_ (.A0(_05523_),
    .A1(_05524_),
    .S(_04817_),
    .X(_05525_));
 sky130_fd_sc_hd__mux2_1 _12340_ (.A0(\rbzero.tex_b0[5] ),
    .A1(\rbzero.tex_b0[4] ),
    .S(_04907_),
    .X(_05526_));
 sky130_fd_sc_hd__mux2_1 _12341_ (.A0(\rbzero.tex_b0[7] ),
    .A1(\rbzero.tex_b0[6] ),
    .S(_04892_),
    .X(_05527_));
 sky130_fd_sc_hd__mux2_1 _12342_ (.A0(_05526_),
    .A1(_05527_),
    .S(_04826_),
    .X(_05528_));
 sky130_fd_sc_hd__mux2_1 _12343_ (.A0(_05525_),
    .A1(_05528_),
    .S(_04918_),
    .X(_05529_));
 sky130_fd_sc_hd__mux2_1 _12344_ (.A0(\rbzero.tex_b0[9] ),
    .A1(\rbzero.tex_b0[8] ),
    .S(_04907_),
    .X(_05530_));
 sky130_fd_sc_hd__or2_1 _12345_ (.A(_04826_),
    .B(_05530_),
    .X(_05531_));
 sky130_fd_sc_hd__mux2_1 _12346_ (.A0(\rbzero.tex_b0[11] ),
    .A1(\rbzero.tex_b0[10] ),
    .S(_04893_),
    .X(_05532_));
 sky130_fd_sc_hd__o21a_1 _12347_ (.A1(_05198_),
    .A2(_05532_),
    .B1(_04939_),
    .X(_05533_));
 sky130_fd_sc_hd__mux2_1 _12348_ (.A0(\rbzero.tex_b0[15] ),
    .A1(\rbzero.tex_b0[14] ),
    .S(_04907_),
    .X(_05534_));
 sky130_fd_sc_hd__mux2_1 _12349_ (.A0(\rbzero.tex_b0[13] ),
    .A1(\rbzero.tex_b0[12] ),
    .S(_04907_),
    .X(_05535_));
 sky130_fd_sc_hd__mux2_1 _12350_ (.A0(_05534_),
    .A1(_05535_),
    .S(_04891_),
    .X(_05536_));
 sky130_fd_sc_hd__a221o_1 _12351_ (.A1(_05531_),
    .A2(_05533_),
    .B1(_05536_),
    .B2(_04952_),
    .C1(_04889_),
    .X(_05537_));
 sky130_fd_sc_hd__o211a_1 _12352_ (.A1(_04812_),
    .A2(_05529_),
    .B1(_05537_),
    .C1(_04886_),
    .X(_05538_));
 sky130_fd_sc_hd__a311o_1 _12353_ (.A1(_04823_),
    .A2(_05514_),
    .A3(_05522_),
    .B1(_05538_),
    .C1(_04832_),
    .X(_05539_));
 sky130_fd_sc_hd__a21o_1 _12354_ (.A1(_05038_),
    .A2(_05372_),
    .B1(_05177_),
    .X(_05540_));
 sky130_fd_sc_hd__nand3_1 _12355_ (.A(_05019_),
    .B(_05371_),
    .C(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hd__o21ba_1 _12356_ (.A1(_05029_),
    .A2(_05541_),
    .B1_N(_05043_),
    .X(_05542_));
 sky130_fd_sc_hd__a31o_1 _12357_ (.A1(_05017_),
    .A2(_05506_),
    .A3(_05539_),
    .B1(_05542_),
    .X(_05543_));
 sky130_fd_sc_hd__mux2_1 _12358_ (.A0(_05472_),
    .A1(_05543_),
    .S(_04899_),
    .X(_05544_));
 sky130_fd_sc_hd__or2_1 _12359_ (.A(_05047_),
    .B(_05544_),
    .X(_05545_));
 sky130_fd_sc_hd__inv_2 _12360_ (.A(_05277_),
    .Y(_05546_));
 sky130_fd_sc_hd__o21a_1 _12361_ (.A1(_05546_),
    .A2(_05290_),
    .B1(_05465_),
    .X(_05547_));
 sky130_fd_sc_hd__or3_1 _12362_ (.A(_04702_),
    .B(_04743_),
    .C(_05547_),
    .X(_05548_));
 sky130_fd_sc_hd__a31o_1 _12363_ (.A1(_05379_),
    .A2(_05545_),
    .A3(_05548_),
    .B1(_04650_),
    .X(_05549_));
 sky130_fd_sc_hd__and2_1 _12364_ (.A(_05051_),
    .B(_05056_),
    .X(_05550_));
 sky130_fd_sc_hd__and3b_4 _12365_ (.A_N(_04661_),
    .B(_05549_),
    .C(_05550_),
    .X(_05551_));
 sky130_fd_sc_hd__mux2_4 _12366_ (.A0(\reg_rgb[22] ),
    .A1(_05551_),
    .S(_05058_),
    .X(_05552_));
 sky130_fd_sc_hd__clkbuf_1 _12367_ (.A(_05552_),
    .X(net66));
 sky130_fd_sc_hd__mux2_1 _12368_ (.A0(\rbzero.color_sky[5] ),
    .A1(\rbzero.color_floor[5] ),
    .S(_04825_),
    .X(_05553_));
 sky130_fd_sc_hd__a21oi_1 _12369_ (.A1(_04818_),
    .A2(_05036_),
    .B1(_05177_),
    .Y(_05554_));
 sky130_fd_sc_hd__or3b_1 _12370_ (.A(_05029_),
    .B(_05554_),
    .C_N(\rbzero.row_render.wall[1] ),
    .X(_05555_));
 sky130_fd_sc_hd__o21ai_1 _12371_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_05186_),
    .B1(_05042_),
    .Y(_05556_));
 sky130_fd_sc_hd__a21o_1 _12372_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_05186_),
    .B1(_05556_),
    .X(_05557_));
 sky130_fd_sc_hd__mux2_1 _12373_ (.A0(\rbzero.tex_b1[41] ),
    .A1(\rbzero.tex_b1[40] ),
    .S(_04931_),
    .X(_05558_));
 sky130_fd_sc_hd__mux2_1 _12374_ (.A0(\rbzero.tex_b1[43] ),
    .A1(\rbzero.tex_b1[42] ),
    .S(_04931_),
    .X(_05559_));
 sky130_fd_sc_hd__mux2_1 _12375_ (.A0(_05558_),
    .A1(_05559_),
    .S(_05190_),
    .X(_05560_));
 sky130_fd_sc_hd__mux2_1 _12376_ (.A0(\rbzero.tex_b1[45] ),
    .A1(\rbzero.tex_b1[44] ),
    .S(_04978_),
    .X(_05561_));
 sky130_fd_sc_hd__mux2_1 _12377_ (.A0(\rbzero.tex_b1[47] ),
    .A1(\rbzero.tex_b1[46] ),
    .S(_04893_),
    .X(_05562_));
 sky130_fd_sc_hd__or2_1 _12378_ (.A(_04981_),
    .B(_05562_),
    .X(_05563_));
 sky130_fd_sc_hd__o211a_1 _12379_ (.A1(_04922_),
    .A2(_05561_),
    .B1(_05563_),
    .C1(_04919_),
    .X(_05564_));
 sky130_fd_sc_hd__a211o_1 _12380_ (.A1(_04937_),
    .A2(_05560_),
    .B1(_05564_),
    .C1(_04967_),
    .X(_05565_));
 sky130_fd_sc_hd__mux2_1 _12381_ (.A0(\rbzero.tex_b1[39] ),
    .A1(\rbzero.tex_b1[38] ),
    .S(_04931_),
    .X(_05566_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(\rbzero.tex_b1[37] ),
    .A1(\rbzero.tex_b1[36] ),
    .S(_04893_),
    .X(_05567_));
 sky130_fd_sc_hd__or2_1 _12383_ (.A(_04826_),
    .B(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__o211a_1 _12384_ (.A1(_05199_),
    .A2(_05566_),
    .B1(_05568_),
    .C1(_04952_),
    .X(_05569_));
 sky130_fd_sc_hd__mux2_1 _12385_ (.A0(\rbzero.tex_b1[33] ),
    .A1(\rbzero.tex_b1[32] ),
    .S(_05009_),
    .X(_05570_));
 sky130_fd_sc_hd__and3_1 _12386_ (.A(\rbzero.tex_b1[35] ),
    .B(_04926_),
    .C(_04928_),
    .X(_05571_));
 sky130_fd_sc_hd__a21o_1 _12387_ (.A1(\rbzero.tex_b1[34] ),
    .A2(_04914_),
    .B1(_04981_),
    .X(_05572_));
 sky130_fd_sc_hd__o221a_1 _12388_ (.A1(_05190_),
    .A2(_05570_),
    .B1(_05571_),
    .B2(_05572_),
    .C1(_04940_),
    .X(_05573_));
 sky130_fd_sc_hd__o31a_1 _12389_ (.A1(_04902_),
    .A2(_05569_),
    .A3(_05573_),
    .B1(_04886_),
    .X(_05574_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(\rbzero.tex_b1[61] ),
    .A1(\rbzero.tex_b1[60] ),
    .S(_04931_),
    .X(_05575_));
 sky130_fd_sc_hd__mux2_1 _12391_ (.A0(\rbzero.tex_b1[63] ),
    .A1(\rbzero.tex_b1[62] ),
    .S(_04931_),
    .X(_05576_));
 sky130_fd_sc_hd__mux2_1 _12392_ (.A0(_05575_),
    .A1(_05576_),
    .S(_05190_),
    .X(_05577_));
 sky130_fd_sc_hd__mux2_1 _12393_ (.A0(\rbzero.tex_b1[57] ),
    .A1(\rbzero.tex_b1[56] ),
    .S(_04931_),
    .X(_05578_));
 sky130_fd_sc_hd__and3_1 _12394_ (.A(\rbzero.tex_b1[59] ),
    .B(_04927_),
    .C(_04929_),
    .X(_05579_));
 sky130_fd_sc_hd__a21o_1 _12395_ (.A1(\rbzero.tex_b1[58] ),
    .A2(_04914_),
    .B1(_04981_),
    .X(_05580_));
 sky130_fd_sc_hd__o221a_1 _12396_ (.A1(_04922_),
    .A2(_05578_),
    .B1(_05579_),
    .B2(_05580_),
    .C1(_04940_),
    .X(_05581_));
 sky130_fd_sc_hd__a211o_1 _12397_ (.A1(_04953_),
    .A2(_05577_),
    .B1(_05581_),
    .C1(_04967_),
    .X(_05582_));
 sky130_fd_sc_hd__mux2_1 _12398_ (.A0(\rbzero.tex_b1[53] ),
    .A1(\rbzero.tex_b1[52] ),
    .S(_04931_),
    .X(_05583_));
 sky130_fd_sc_hd__mux2_1 _12399_ (.A0(\rbzero.tex_b1[55] ),
    .A1(\rbzero.tex_b1[54] ),
    .S(_04893_),
    .X(_05584_));
 sky130_fd_sc_hd__or2_1 _12400_ (.A(_05198_),
    .B(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__o211a_1 _12401_ (.A1(_05190_),
    .A2(_05583_),
    .B1(_05585_),
    .C1(_04952_),
    .X(_05586_));
 sky130_fd_sc_hd__mux2_1 _12402_ (.A0(\rbzero.tex_b1[49] ),
    .A1(\rbzero.tex_b1[48] ),
    .S(_05314_),
    .X(_05587_));
 sky130_fd_sc_hd__mux2_1 _12403_ (.A0(\rbzero.tex_b1[51] ),
    .A1(\rbzero.tex_b1[50] ),
    .S(_04893_),
    .X(_05588_));
 sky130_fd_sc_hd__or2_1 _12404_ (.A(_05198_),
    .B(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__o211a_1 _12405_ (.A1(_04922_),
    .A2(_05587_),
    .B1(_05589_),
    .C1(_04940_),
    .X(_05590_));
 sky130_fd_sc_hd__o31a_1 _12406_ (.A1(_04902_),
    .A2(_05586_),
    .A3(_05590_),
    .B1(_04823_),
    .X(_05591_));
 sky130_fd_sc_hd__a221o_1 _12407_ (.A1(_05565_),
    .A2(_05574_),
    .B1(_05582_),
    .B2(_05591_),
    .C1(_04810_),
    .X(_05592_));
 sky130_fd_sc_hd__mux2_1 _12408_ (.A0(\rbzero.tex_b1[9] ),
    .A1(\rbzero.tex_b1[8] ),
    .S(_04978_),
    .X(_05593_));
 sky130_fd_sc_hd__mux2_1 _12409_ (.A0(\rbzero.tex_b1[11] ),
    .A1(\rbzero.tex_b1[10] ),
    .S(_05314_),
    .X(_05594_));
 sky130_fd_sc_hd__mux2_1 _12410_ (.A0(_05593_),
    .A1(_05594_),
    .S(_05190_),
    .X(_05595_));
 sky130_fd_sc_hd__mux2_1 _12411_ (.A0(\rbzero.tex_b1[13] ),
    .A1(\rbzero.tex_b1[12] ),
    .S(_04978_),
    .X(_05596_));
 sky130_fd_sc_hd__mux2_1 _12412_ (.A0(\rbzero.tex_b1[15] ),
    .A1(\rbzero.tex_b1[14] ),
    .S(_04913_),
    .X(_05597_));
 sky130_fd_sc_hd__or2_1 _12413_ (.A(_04981_),
    .B(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__o211a_1 _12414_ (.A1(_04944_),
    .A2(_05596_),
    .B1(_05598_),
    .C1(_04919_),
    .X(_05599_));
 sky130_fd_sc_hd__a211o_1 _12415_ (.A1(_04937_),
    .A2(_05595_),
    .B1(_05599_),
    .C1(_04967_),
    .X(_05600_));
 sky130_fd_sc_hd__mux2_1 _12416_ (.A0(\rbzero.tex_b1[5] ),
    .A1(\rbzero.tex_b1[4] ),
    .S(_05314_),
    .X(_05601_));
 sky130_fd_sc_hd__mux2_1 _12417_ (.A0(\rbzero.tex_b1[7] ),
    .A1(\rbzero.tex_b1[6] ),
    .S(_05314_),
    .X(_05602_));
 sky130_fd_sc_hd__mux2_1 _12418_ (.A0(_05601_),
    .A1(_05602_),
    .S(_05190_),
    .X(_05603_));
 sky130_fd_sc_hd__mux2_1 _12419_ (.A0(\rbzero.tex_b1[1] ),
    .A1(\rbzero.tex_b1[0] ),
    .S(_05314_),
    .X(_05604_));
 sky130_fd_sc_hd__and3_1 _12420_ (.A(\rbzero.tex_b1[3] ),
    .B(_04927_),
    .C(_04929_),
    .X(_05605_));
 sky130_fd_sc_hd__a21o_1 _12421_ (.A1(\rbzero.tex_b1[2] ),
    .A2(_04909_),
    .B1(_04981_),
    .X(_05606_));
 sky130_fd_sc_hd__o221a_1 _12422_ (.A1(_04922_),
    .A2(_05604_),
    .B1(_05605_),
    .B2(_05606_),
    .C1(_04940_),
    .X(_05607_));
 sky130_fd_sc_hd__a211o_1 _12423_ (.A1(_04953_),
    .A2(_05603_),
    .B1(_05607_),
    .C1(_04902_),
    .X(_05608_));
 sky130_fd_sc_hd__mux2_1 _12424_ (.A0(\rbzero.tex_b1[29] ),
    .A1(\rbzero.tex_b1[28] ),
    .S(_04913_),
    .X(_05609_));
 sky130_fd_sc_hd__mux2_1 _12425_ (.A0(\rbzero.tex_b1[31] ),
    .A1(\rbzero.tex_b1[30] ),
    .S(_04913_),
    .X(_05610_));
 sky130_fd_sc_hd__mux2_1 _12426_ (.A0(_05609_),
    .A1(_05610_),
    .S(_04826_),
    .X(_05611_));
 sky130_fd_sc_hd__mux2_1 _12427_ (.A0(\rbzero.tex_b1[25] ),
    .A1(\rbzero.tex_b1[24] ),
    .S(_04893_),
    .X(_05612_));
 sky130_fd_sc_hd__and3_1 _12428_ (.A(\rbzero.tex_b1[27] ),
    .B(_04926_),
    .C(_04928_),
    .X(_05613_));
 sky130_fd_sc_hd__a21o_1 _12429_ (.A1(\rbzero.tex_b1[26] ),
    .A2(_04908_),
    .B1(_04817_),
    .X(_05614_));
 sky130_fd_sc_hd__o221a_1 _12430_ (.A1(_04827_),
    .A2(_05612_),
    .B1(_05613_),
    .B2(_05614_),
    .C1(_04939_),
    .X(_05615_));
 sky130_fd_sc_hd__a211o_1 _12431_ (.A1(_04919_),
    .A2(_05611_),
    .B1(_05615_),
    .C1(_04889_),
    .X(_05616_));
 sky130_fd_sc_hd__mux2_1 _12432_ (.A0(\rbzero.tex_b1[17] ),
    .A1(\rbzero.tex_b1[16] ),
    .S(_04913_),
    .X(_05617_));
 sky130_fd_sc_hd__mux2_1 _12433_ (.A0(\rbzero.tex_b1[19] ),
    .A1(\rbzero.tex_b1[18] ),
    .S(_04893_),
    .X(_05618_));
 sky130_fd_sc_hd__mux2_1 _12434_ (.A0(_05617_),
    .A1(_05618_),
    .S(_04826_),
    .X(_05619_));
 sky130_fd_sc_hd__mux2_1 _12435_ (.A0(\rbzero.tex_b1[21] ),
    .A1(\rbzero.tex_b1[20] ),
    .S(_04913_),
    .X(_05620_));
 sky130_fd_sc_hd__mux2_1 _12436_ (.A0(\rbzero.tex_b1[23] ),
    .A1(\rbzero.tex_b1[22] ),
    .S(_04892_),
    .X(_05621_));
 sky130_fd_sc_hd__or2_1 _12437_ (.A(_04817_),
    .B(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__o211a_1 _12438_ (.A1(_04827_),
    .A2(_05620_),
    .B1(_05622_),
    .C1(_04918_),
    .X(_05623_));
 sky130_fd_sc_hd__a211o_1 _12439_ (.A1(_04940_),
    .A2(_05619_),
    .B1(_05623_),
    .C1(_04812_),
    .X(_05624_));
 sky130_fd_sc_hd__a31o_1 _12440_ (.A1(_04823_),
    .A2(_05616_),
    .A3(_05624_),
    .B1(_04832_),
    .X(_05625_));
 sky130_fd_sc_hd__a31o_1 _12441_ (.A1(_04887_),
    .A2(_05600_),
    .A3(_05608_),
    .B1(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__a21oi_2 _12442_ (.A1(_05592_),
    .A2(_05626_),
    .B1(_05263_),
    .Y(_05627_));
 sky130_fd_sc_hd__a31o_1 _12443_ (.A1(_05263_),
    .A2(_05555_),
    .A3(_05557_),
    .B1(_05627_),
    .X(_05628_));
 sky130_fd_sc_hd__nand2_1 _12444_ (.A(_04900_),
    .B(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__o211a_1 _12445_ (.A1(_04900_),
    .A2(_05553_),
    .B1(_05629_),
    .C1(_04702_),
    .X(_05630_));
 sky130_fd_sc_hd__a311o_1 _12446_ (.A1(_05047_),
    .A2(_04744_),
    .A3(_05547_),
    .B1(_05630_),
    .C1(_04650_),
    .X(_05631_));
 sky130_fd_sc_hd__and3b_4 _12447_ (.A_N(_05176_),
    .B(_05550_),
    .C(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__mux2_4 _12448_ (.A0(\reg_rgb[23] ),
    .A1(_05632_),
    .S(_05058_),
    .X(_05633_));
 sky130_fd_sc_hd__clkbuf_1 _12449_ (.A(_05633_),
    .X(net67));
 sky130_fd_sc_hd__mux2_2 _12450_ (.A0(reg_vsync),
    .A1(_04431_),
    .S(_05058_),
    .X(_05634_));
 sky130_fd_sc_hd__clkbuf_1 _12451_ (.A(_05634_),
    .X(net74));
 sky130_fd_sc_hd__clkinv_2 _12452_ (.A(\rbzero.hsync ),
    .Y(_05635_));
 sky130_fd_sc_hd__mux2_2 _12453_ (.A0(reg_hsync),
    .A1(_05635_),
    .S(_05058_),
    .X(_05636_));
 sky130_fd_sc_hd__clkbuf_1 _12454_ (.A(_05636_),
    .X(net62));
 sky130_fd_sc_hd__nor2_1 _12455_ (.A(net5),
    .B(net4),
    .Y(_05637_));
 sky130_fd_sc_hd__nor2_2 _12456_ (.A(net7),
    .B(net6),
    .Y(_05638_));
 sky130_fd_sc_hd__nand2_1 _12457_ (.A(_05637_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__buf_2 _12458_ (.A(net6),
    .X(_05640_));
 sky130_fd_sc_hd__a21o_1 _12459_ (.A1(net5),
    .A2(_05640_),
    .B1(net7),
    .X(_05641_));
 sky130_fd_sc_hd__nand2_1 _12460_ (.A(net8),
    .B(_05641_),
    .Y(_05642_));
 sky130_fd_sc_hd__inv_2 _12461_ (.A(net5),
    .Y(_05643_));
 sky130_fd_sc_hd__buf_2 _12462_ (.A(_04653_),
    .X(_05644_));
 sky130_fd_sc_hd__buf_2 _12463_ (.A(_04648_),
    .X(_05645_));
 sky130_fd_sc_hd__clkbuf_4 _12464_ (.A(net4),
    .X(_05646_));
 sky130_fd_sc_hd__mux4_1 _12465_ (.A0(_04687_),
    .A1(_05644_),
    .A2(_05645_),
    .A3(_04642_),
    .S0(_05646_),
    .S1(_05640_),
    .X(_05647_));
 sky130_fd_sc_hd__buf_2 _12466_ (.A(_04651_),
    .X(_05648_));
 sky130_fd_sc_hd__mux2_1 _12467_ (.A0(_05648_),
    .A1(_04657_),
    .S(_05646_),
    .X(_05649_));
 sky130_fd_sc_hd__clkbuf_4 _12468_ (.A(\gpout0.vpos[0] ),
    .X(_05650_));
 sky130_fd_sc_hd__buf_2 _12469_ (.A(\gpout0.vpos[1] ),
    .X(_05651_));
 sky130_fd_sc_hd__clkbuf_4 _12470_ (.A(\gpout0.vpos[8] ),
    .X(_05652_));
 sky130_fd_sc_hd__buf_2 _12471_ (.A(\gpout0.vpos[9] ),
    .X(_05653_));
 sky130_fd_sc_hd__mux4_1 _12472_ (.A0(_05650_),
    .A1(_05651_),
    .A2(_05652_),
    .A3(_05653_),
    .S0(_05646_),
    .S1(net7),
    .X(_05654_));
 sky130_fd_sc_hd__or2b_1 _12473_ (.A(_05654_),
    .B_N(_05640_),
    .X(_05655_));
 sky130_fd_sc_hd__o211a_1 _12474_ (.A1(_05640_),
    .A2(_05649_),
    .B1(_05655_),
    .C1(net5),
    .X(_05656_));
 sky130_fd_sc_hd__a21oi_1 _12475_ (.A1(_05643_),
    .A2(_05647_),
    .B1(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__inv_2 _12476_ (.A(net4),
    .Y(_05658_));
 sky130_fd_sc_hd__nor2_1 _12477_ (.A(net5),
    .B(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__a22oi_1 _12478_ (.A1(_05055_),
    .A2(_05637_),
    .B1(_05659_),
    .B2(net71),
    .Y(_05660_));
 sky130_fd_sc_hd__inv_2 _12479_ (.A(net7),
    .Y(_05661_));
 sky130_fd_sc_hd__nand2_1 _12480_ (.A(_05661_),
    .B(_05640_),
    .Y(_05662_));
 sky130_fd_sc_hd__nor2_1 _12481_ (.A(_05643_),
    .B(_05658_),
    .Y(_05663_));
 sky130_fd_sc_hd__nor2_1 _12482_ (.A(_05643_),
    .B(_05646_),
    .Y(_05664_));
 sky130_fd_sc_hd__nor2_1 _12483_ (.A(net9),
    .B(net8),
    .Y(_05665_));
 sky130_fd_sc_hd__and3_1 _12484_ (.A(net54),
    .B(_05663_),
    .C(_05665_),
    .X(_05666_));
 sky130_fd_sc_hd__a221o_1 _12485_ (.A1(net49),
    .A2(_05664_),
    .B1(_05663_),
    .B2(net50),
    .C1(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__a22o_1 _12486_ (.A1(net51),
    .A2(_05637_),
    .B1(_05659_),
    .B2(net40),
    .X(_05668_));
 sky130_fd_sc_hd__a221o_1 _12487_ (.A1(net41),
    .A2(_05664_),
    .B1(_05663_),
    .B2(_05263_),
    .C1(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__and3b_1 _12488_ (.A_N(net6),
    .B(_05669_),
    .C(net7),
    .X(_05670_));
 sky130_fd_sc_hd__a31o_1 _12489_ (.A1(net43),
    .A2(_05637_),
    .A3(_05638_),
    .B1(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__a31o_1 _12490_ (.A1(_05661_),
    .A2(_05640_),
    .A3(_05667_),
    .B1(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__a31o_1 _12491_ (.A1(net46),
    .A2(_05659_),
    .A3(_05638_),
    .B1(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__and3_1 _12492_ (.A(net44),
    .B(_05664_),
    .C(_05638_),
    .X(_05674_));
 sky130_fd_sc_hd__a311o_1 _12493_ (.A1(_05053_),
    .A2(_05638_),
    .A3(_05663_),
    .B1(_05673_),
    .C1(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__o21ba_1 _12494_ (.A1(_05660_),
    .A2(_05662_),
    .B1_N(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__o22ai_1 _12495_ (.A1(_05642_),
    .A2(_05657_),
    .B1(_05676_),
    .B2(net8),
    .Y(_05677_));
 sky130_fd_sc_hd__a21o_1 _12496_ (.A1(net7),
    .A2(_05640_),
    .B1(net8),
    .X(_05678_));
 sky130_fd_sc_hd__mux4_1 _12497_ (.A0(_04589_),
    .A1(_04704_),
    .A2(_04419_),
    .A3(_03973_),
    .S0(_05646_),
    .S1(net5),
    .X(_05679_));
 sky130_fd_sc_hd__mux4_1 _12498_ (.A0(_03969_),
    .A1(\gpout0.hpos[1] ),
    .A2(_04452_),
    .A3(_04628_),
    .S0(_05646_),
    .S1(net5),
    .X(_05680_));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(_03975_),
    .A1(_04420_),
    .S(_05646_),
    .X(_05681_));
 sky130_fd_sc_hd__mux2_1 _12500_ (.A0(_05680_),
    .A1(_05681_),
    .S(_05661_),
    .X(_05682_));
 sky130_fd_sc_hd__mux2_1 _12501_ (.A0(_05679_),
    .A1(_05682_),
    .S(_05640_),
    .X(_05683_));
 sky130_fd_sc_hd__a22o_1 _12502_ (.A1(net52),
    .A2(_05637_),
    .B1(_05664_),
    .B2(net55),
    .X(_05684_));
 sky130_fd_sc_hd__a21oi_1 _12503_ (.A1(net53),
    .A2(_05659_),
    .B1(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__nor2_1 _12504_ (.A(_05662_),
    .B(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__o211a_1 _12505_ (.A1(_05658_),
    .A2(_04052_),
    .B1(_05638_),
    .C1(_05643_),
    .X(_05687_));
 sky130_fd_sc_hd__and3_2 _12506_ (.A(clknet_3_3_0_i_clk),
    .B(_05664_),
    .C(_05638_),
    .X(_05688_));
 sky130_fd_sc_hd__a31o_2 _12507_ (.A1(\gpout0.clk_div[1] ),
    .A2(_05638_),
    .A3(_05663_),
    .B1(_05688_),
    .X(_05689_));
 sky130_fd_sc_hd__o31a_2 _12508_ (.A1(_05686_),
    .A2(_05687_),
    .A3(_05689_),
    .B1(_05665_),
    .X(_05690_));
 sky130_fd_sc_hd__a41o_2 _12509_ (.A1(net9),
    .A2(_05642_),
    .A3(_05678_),
    .A4(_05683_),
    .B1(_05690_),
    .X(_05691_));
 sky130_fd_sc_hd__a31o_2 _12510_ (.A1(_05661_),
    .A2(_05640_),
    .A3(_05666_),
    .B1(_05691_),
    .X(_05692_));
 sky130_fd_sc_hd__or2_1 _12511_ (.A(_05646_),
    .B(_05057_),
    .X(_05693_));
 sky130_fd_sc_hd__nor2_1 _12512_ (.A(_05661_),
    .B(net8),
    .Y(_05694_));
 sky130_fd_sc_hd__nand2_1 _12513_ (.A(_05646_),
    .B(_05297_),
    .Y(_05695_));
 sky130_fd_sc_hd__mux4_1 _12514_ (.A0(_05382_),
    .A1(_05470_),
    .A2(_05551_),
    .A3(_05632_),
    .S0(_05646_),
    .S1(net7),
    .X(_05696_));
 sky130_fd_sc_hd__a32o_1 _12515_ (.A1(_05693_),
    .A2(_05694_),
    .A3(_05695_),
    .B1(_05696_),
    .B2(net8),
    .X(_05697_));
 sky130_fd_sc_hd__and4b_1 _12516_ (.A_N(net9),
    .B(_05697_),
    .C(net5),
    .D(_05640_),
    .X(_05698_));
 sky130_fd_sc_hd__a211o_2 _12517_ (.A1(net9),
    .A2(_05677_),
    .B1(_05692_),
    .C1(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__o41a_2 _12518_ (.A1(net9),
    .A2(net8),
    .A3(_05382_),
    .A4(_05639_),
    .B1(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__mux2_2 _12519_ (.A0(\reg_gpout[0] ),
    .A1(clknet_1_1__leaf__05700_),
    .S(_05058_),
    .X(_05701_));
 sky130_fd_sc_hd__buf_1 _12520_ (.A(_05701_),
    .X(net56));
 sky130_fd_sc_hd__inv_2 _12521_ (.A(net11),
    .Y(_05702_));
 sky130_fd_sc_hd__inv_2 _12522_ (.A(net12),
    .Y(_05703_));
 sky130_fd_sc_hd__buf_2 _12523_ (.A(net10),
    .X(_05704_));
 sky130_fd_sc_hd__mux4_1 _12524_ (.A0(_05382_),
    .A1(_05470_),
    .A2(_05551_),
    .A3(_05632_),
    .S0(_05704_),
    .S1(net13),
    .X(_05705_));
 sky130_fd_sc_hd__nand2_1 _12525_ (.A(_05704_),
    .B(_05297_),
    .Y(_05706_));
 sky130_fd_sc_hd__inv_2 _12526_ (.A(net14),
    .Y(_05707_));
 sky130_fd_sc_hd__o2111a_1 _12527_ (.A1(_05704_),
    .A2(_05057_),
    .B1(_05706_),
    .C1(net13),
    .D1(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__a21oi_1 _12528_ (.A1(net14),
    .A2(_05705_),
    .B1(_05708_),
    .Y(_05709_));
 sky130_fd_sc_hd__or4_1 _12529_ (.A(_05702_),
    .B(_05703_),
    .C(net15),
    .D(_05709_),
    .X(_05710_));
 sky130_fd_sc_hd__clkbuf_8 _12530_ (.A(net54),
    .X(_05711_));
 sky130_fd_sc_hd__and2_1 _12531_ (.A(net11),
    .B(_05704_),
    .X(_05712_));
 sky130_fd_sc_hd__nor2_1 _12532_ (.A(net14),
    .B(net15),
    .Y(_05713_));
 sky130_fd_sc_hd__and3_1 _12533_ (.A(_05711_),
    .B(_05712_),
    .C(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__nor2_2 _12534_ (.A(_05702_),
    .B(_05704_),
    .Y(_05715_));
 sky130_fd_sc_hd__a22o_1 _12535_ (.A1(net50),
    .A2(_05712_),
    .B1(_05715_),
    .B2(net49),
    .X(_05716_));
 sky130_fd_sc_hd__inv_2 _12536_ (.A(net13),
    .Y(_05717_));
 sky130_fd_sc_hd__o21a_1 _12537_ (.A1(_05714_),
    .A2(_05716_),
    .B1(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__nor2_2 _12538_ (.A(net11),
    .B(net10),
    .Y(_05719_));
 sky130_fd_sc_hd__and2_1 _12539_ (.A(_05702_),
    .B(_05704_),
    .X(_05720_));
 sky130_fd_sc_hd__nor2_1 _12540_ (.A(net13),
    .B(net12),
    .Y(_05721_));
 sky130_fd_sc_hd__inv_2 _12541_ (.A(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__a221o_1 _12542_ (.A1(net43),
    .A2(_05719_),
    .B1(_05720_),
    .B2(net46),
    .C1(_05722_),
    .X(_05723_));
 sky130_fd_sc_hd__a22o_1 _12543_ (.A1(net40),
    .A2(_05720_),
    .B1(_05715_),
    .B2(net41),
    .X(_05724_));
 sky130_fd_sc_hd__a221o_1 _12544_ (.A1(net51),
    .A2(_05719_),
    .B1(_05712_),
    .B2(_05263_),
    .C1(_05717_),
    .X(_05725_));
 sky130_fd_sc_hd__nor2_1 _12545_ (.A(net13),
    .B(_05703_),
    .Y(_05726_));
 sky130_fd_sc_hd__a31o_1 _12546_ (.A1(_05711_),
    .A2(_05726_),
    .A3(_05712_),
    .B1(net15),
    .X(_05727_));
 sky130_fd_sc_hd__o21a_1 _12547_ (.A1(_05724_),
    .A2(_05725_),
    .B1(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__o2111a_1 _12548_ (.A1(_05703_),
    .A2(_05718_),
    .B1(_05723_),
    .C1(_05728_),
    .D1(_05707_),
    .X(_05729_));
 sky130_fd_sc_hd__or2b_1 _12549_ (.A(\gpout0.vpos[1] ),
    .B_N(net10),
    .X(_05730_));
 sky130_fd_sc_hd__o2111a_1 _12550_ (.A1(_05650_),
    .A2(_05704_),
    .B1(net12),
    .C1(_05730_),
    .D1(net11),
    .X(_05731_));
 sky130_fd_sc_hd__nand2_1 _12551_ (.A(_05702_),
    .B(net10),
    .Y(_05732_));
 sky130_fd_sc_hd__mux2_1 _12552_ (.A0(_04419_),
    .A1(_03973_),
    .S(net10),
    .X(_05733_));
 sky130_fd_sc_hd__or2_1 _12553_ (.A(_05702_),
    .B(_05733_),
    .X(_05734_));
 sky130_fd_sc_hd__nand2_1 _12554_ (.A(_04414_),
    .B(_05719_),
    .Y(_05735_));
 sky130_fd_sc_hd__o2111a_1 _12555_ (.A1(_04704_),
    .A2(_05732_),
    .B1(_05734_),
    .C1(_05703_),
    .D1(_05735_),
    .X(_05736_));
 sky130_fd_sc_hd__nor2_1 _12556_ (.A(_03975_),
    .B(_05704_),
    .Y(_05737_));
 sky130_fd_sc_hd__a2111oi_1 _12557_ (.A1(_03976_),
    .A2(_05704_),
    .B1(_05703_),
    .C1(_05737_),
    .D1(net11),
    .Y(_05738_));
 sky130_fd_sc_hd__o31a_1 _12558_ (.A1(_05731_),
    .A2(_05736_),
    .A3(_05738_),
    .B1(_05717_),
    .X(_05739_));
 sky130_fd_sc_hd__mux4_1 _12559_ (.A0(_04651_),
    .A1(_04657_),
    .A2(_05652_),
    .A3(_05653_),
    .S0(net10),
    .S1(net12),
    .X(_05740_));
 sky130_fd_sc_hd__mux4_1 _12560_ (.A0(_04687_),
    .A1(_04653_),
    .A2(_05645_),
    .A3(_04642_),
    .S0(net10),
    .S1(net12),
    .X(_05741_));
 sky130_fd_sc_hd__or2_1 _12561_ (.A(net11),
    .B(_05741_),
    .X(_05742_));
 sky130_fd_sc_hd__o211a_1 _12562_ (.A1(_05702_),
    .A2(_05740_),
    .B1(_05742_),
    .C1(net13),
    .X(_05743_));
 sky130_fd_sc_hd__or3_1 _12563_ (.A(_05707_),
    .B(_05739_),
    .C(_05743_),
    .X(_05744_));
 sky130_fd_sc_hd__a22o_1 _12564_ (.A1(_05055_),
    .A2(_05719_),
    .B1(_05720_),
    .B2(net71),
    .X(_05745_));
 sky130_fd_sc_hd__a22o_1 _12565_ (.A1(_05053_),
    .A2(_05712_),
    .B1(_05715_),
    .B2(net44),
    .X(_05746_));
 sky130_fd_sc_hd__a221o_1 _12566_ (.A1(_05726_),
    .A2(_05745_),
    .B1(_05721_),
    .B2(_05746_),
    .C1(net14),
    .X(_05747_));
 sky130_fd_sc_hd__a2111oi_1 _12567_ (.A1(_04454_),
    .A2(_05719_),
    .B1(net14),
    .C1(_05703_),
    .D1(_05717_),
    .Y(_05748_));
 sky130_fd_sc_hd__nand2_1 _12568_ (.A(net11),
    .B(_05704_),
    .Y(_05749_));
 sky130_fd_sc_hd__nand2_1 _12569_ (.A(_04446_),
    .B(_05715_),
    .Y(_05750_));
 sky130_fd_sc_hd__o221a_1 _12570_ (.A1(_04575_),
    .A2(_05732_),
    .B1(_05749_),
    .B2(_04628_),
    .C1(_05750_),
    .X(_05751_));
 sky130_fd_sc_hd__a22o_1 _12571_ (.A1(_05744_),
    .A2(_05747_),
    .B1(_05748_),
    .B2(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__and2_1 _12572_ (.A(net52),
    .B(_05719_),
    .X(_05753_));
 sky130_fd_sc_hd__a221o_1 _12573_ (.A1(net53),
    .A2(_05720_),
    .B1(_05715_),
    .B2(net55),
    .C1(_05753_),
    .X(_05754_));
 sky130_fd_sc_hd__inv_2 _12574_ (.A(_05715_),
    .Y(_05755_));
 sky130_fd_sc_hd__o221a_2 _12575_ (.A1(\gpout1.clk_div[1] ),
    .A2(_05749_),
    .B1(_05755_),
    .B2(clknet_1_0__leaf__04634_),
    .C1(_05721_),
    .X(_05756_));
 sky130_fd_sc_hd__a21o_2 _12576_ (.A1(_05726_),
    .A2(_05754_),
    .B1(_05756_),
    .X(_05757_));
 sky130_fd_sc_hd__a22o_2 _12577_ (.A1(net15),
    .A2(_05752_),
    .B1(_05713_),
    .B2(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__nor2_2 _12578_ (.A(_05729_),
    .B(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__and4b_1 _12579_ (.A_N(_05470_),
    .B(_05719_),
    .C(_05721_),
    .D(_05713_),
    .X(_05760_));
 sky130_fd_sc_hd__a21oi_2 _12580_ (.A1(_05710_),
    .A2(_05759_),
    .B1(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__mux2_2 _12581_ (.A0(\reg_gpout[1] ),
    .A1(clknet_1_1__leaf__05761_),
    .S(_05058_),
    .X(_05762_));
 sky130_fd_sc_hd__buf_1 _12582_ (.A(_05762_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 _12583_ (.A(net16),
    .X(_05763_));
 sky130_fd_sc_hd__or2_1 _12584_ (.A(_05763_),
    .B(_05057_),
    .X(_05764_));
 sky130_fd_sc_hd__inv_2 _12585_ (.A(net19),
    .Y(_05765_));
 sky130_fd_sc_hd__nor2_1 _12586_ (.A(_05765_),
    .B(net20),
    .Y(_05766_));
 sky130_fd_sc_hd__nand2_1 _12587_ (.A(_05763_),
    .B(_05297_),
    .Y(_05767_));
 sky130_fd_sc_hd__mux4_1 _12588_ (.A0(_05382_),
    .A1(_05470_),
    .A2(_05551_),
    .A3(_05632_),
    .S0(_05763_),
    .S1(net19),
    .X(_05768_));
 sky130_fd_sc_hd__a32o_1 _12589_ (.A1(_05764_),
    .A2(_05766_),
    .A3(_05767_),
    .B1(_05768_),
    .B2(net20),
    .X(_05769_));
 sky130_fd_sc_hd__buf_2 _12590_ (.A(net18),
    .X(_05770_));
 sky130_fd_sc_hd__and4b_1 _12591_ (.A_N(net21),
    .B(_05769_),
    .C(net17),
    .D(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__a21oi_1 _12592_ (.A1(net17),
    .A2(_05770_),
    .B1(net19),
    .Y(_05772_));
 sky130_fd_sc_hd__a22o_1 _12593_ (.A1(_05770_),
    .A2(_05766_),
    .B1(_05772_),
    .B2(net20),
    .X(_05773_));
 sky130_fd_sc_hd__mux4_1 _12594_ (.A0(_04589_),
    .A1(_04704_),
    .A2(_04419_),
    .A3(_03973_),
    .S0(_05763_),
    .S1(net17),
    .X(_05774_));
 sky130_fd_sc_hd__mux4_1 _12595_ (.A0(_03969_),
    .A1(\gpout0.hpos[1] ),
    .A2(_04452_),
    .A3(_04628_),
    .S0(net16),
    .S1(net17),
    .X(_05775_));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(_03975_),
    .A1(_04420_),
    .S(_05763_),
    .X(_05776_));
 sky130_fd_sc_hd__mux2_1 _12597_ (.A0(_05775_),
    .A1(_05776_),
    .S(_05765_),
    .X(_05777_));
 sky130_fd_sc_hd__mux2_1 _12598_ (.A0(_05774_),
    .A1(_05777_),
    .S(_05770_),
    .X(_05778_));
 sky130_fd_sc_hd__and3_1 _12599_ (.A(net21),
    .B(_05773_),
    .C(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__inv_2 _12600_ (.A(net17),
    .Y(_05780_));
 sky130_fd_sc_hd__mux4_1 _12601_ (.A0(_04687_),
    .A1(_05644_),
    .A2(_05645_),
    .A3(_04642_),
    .S0(_05763_),
    .S1(_05770_),
    .X(_05781_));
 sky130_fd_sc_hd__inv_2 _12602_ (.A(_05770_),
    .Y(_05782_));
 sky130_fd_sc_hd__mux4_1 _12603_ (.A0(_05650_),
    .A1(_05651_),
    .A2(_05652_),
    .A3(_05653_),
    .S0(net16),
    .S1(net19),
    .X(_05783_));
 sky130_fd_sc_hd__or2_1 _12604_ (.A(_05782_),
    .B(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__mux2_1 _12605_ (.A0(_05648_),
    .A1(_04657_),
    .S(_05763_),
    .X(_05785_));
 sky130_fd_sc_hd__o21a_1 _12606_ (.A1(_05770_),
    .A2(_05785_),
    .B1(net17),
    .X(_05786_));
 sky130_fd_sc_hd__a22o_1 _12607_ (.A1(_05780_),
    .A2(_05781_),
    .B1(_05784_),
    .B2(_05786_),
    .X(_05787_));
 sky130_fd_sc_hd__and4b_1 _12608_ (.A_N(_05772_),
    .B(_05787_),
    .C(net21),
    .D(net20),
    .X(_05788_));
 sky130_fd_sc_hd__mux4_1 _12609_ (.A0(net51),
    .A1(net41),
    .A2(net40),
    .A3(_05263_),
    .S0(net17),
    .S1(_05763_),
    .X(_05789_));
 sky130_fd_sc_hd__nor2_1 _12610_ (.A(net19),
    .B(net18),
    .Y(_05790_));
 sky130_fd_sc_hd__nor2_1 _12611_ (.A(_05780_),
    .B(_05763_),
    .Y(_05791_));
 sky130_fd_sc_hd__nand2_1 _12612_ (.A(net17),
    .B(_05763_),
    .Y(_05792_));
 sky130_fd_sc_hd__nor2_1 _12613_ (.A(net21),
    .B(net20),
    .Y(_05793_));
 sky130_fd_sc_hd__a21oi_1 _12614_ (.A1(_05711_),
    .A2(_05793_),
    .B1(net50),
    .Y(_05794_));
 sky130_fd_sc_hd__o2bb2a_1 _12615_ (.A1_N(net49),
    .A2_N(_05791_),
    .B1(_05792_),
    .B2(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__nor2_1 _12616_ (.A(net19),
    .B(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__a211o_1 _12617_ (.A1(_05782_),
    .A2(_05789_),
    .B1(_05790_),
    .C1(_05796_),
    .X(_05797_));
 sky130_fd_sc_hd__and3b_1 _12618_ (.A_N(_05792_),
    .B(_05765_),
    .C(_05770_),
    .X(_05798_));
 sky130_fd_sc_hd__and2b_1 _12619_ (.A_N(net20),
    .B(net21),
    .X(_05799_));
 sky130_fd_sc_hd__a31o_1 _12620_ (.A1(_05711_),
    .A2(_05793_),
    .A3(_05798_),
    .B1(_05799_),
    .X(_05800_));
 sky130_fd_sc_hd__inv_2 _12621_ (.A(net16),
    .Y(_05801_));
 sky130_fd_sc_hd__nor2_1 _12622_ (.A(net17),
    .B(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__nor2_1 _12623_ (.A(net17),
    .B(net16),
    .Y(_05803_));
 sky130_fd_sc_hd__or2_1 _12624_ (.A(net19),
    .B(net18),
    .X(_05804_));
 sky130_fd_sc_hd__a221o_1 _12625_ (.A1(net46),
    .A2(_05802_),
    .B1(_05803_),
    .B2(net43),
    .C1(_05804_),
    .X(_05805_));
 sky130_fd_sc_hd__and2_1 _12626_ (.A(net52),
    .B(_05803_),
    .X(_05806_));
 sky130_fd_sc_hd__a221o_1 _12627_ (.A1(net55),
    .A2(_05791_),
    .B1(_05802_),
    .B2(net53),
    .C1(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__nor2_1 _12628_ (.A(_05792_),
    .B(_05804_),
    .Y(_05808_));
 sky130_fd_sc_hd__o211a_1 _12629_ (.A1(net47),
    .A2(_05801_),
    .B1(_05790_),
    .C1(_05780_),
    .X(_05809_));
 sky130_fd_sc_hd__and3_2 _12630_ (.A(clknet_leaf_40_i_clk),
    .B(_05791_),
    .C(_05790_),
    .X(_05810_));
 sky130_fd_sc_hd__a211o_2 _12631_ (.A1(\gpout2.clk_div[1] ),
    .A2(_05808_),
    .B1(_05809_),
    .C1(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__a31o_2 _12632_ (.A1(_05765_),
    .A2(_05770_),
    .A3(_05807_),
    .B1(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__a32o_2 _12633_ (.A1(_05797_),
    .A2(_05800_),
    .A3(_05805_),
    .B1(_05812_),
    .B2(_05793_),
    .X(_05813_));
 sky130_fd_sc_hd__a22o_1 _12634_ (.A1(net71),
    .A2(_05802_),
    .B1(_05803_),
    .B2(_05055_),
    .X(_05814_));
 sky130_fd_sc_hd__a32o_1 _12635_ (.A1(net44),
    .A2(_05791_),
    .A3(_05790_),
    .B1(_05808_),
    .B2(_05053_),
    .X(_05815_));
 sky130_fd_sc_hd__a31o_1 _12636_ (.A1(_05765_),
    .A2(_05770_),
    .A3(_05814_),
    .B1(_05815_),
    .X(_05816_));
 sky130_fd_sc_hd__nand2_1 _12637_ (.A(_05799_),
    .B(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__or4b_2 _12638_ (.A(_05779_),
    .B(_05788_),
    .C(_05813_),
    .D_N(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__nand3_1 _12639_ (.A(_05793_),
    .B(_05803_),
    .C(_05790_),
    .Y(_05819_));
 sky130_fd_sc_hd__o22a_2 _12640_ (.A1(_05771_),
    .A2(_05818_),
    .B1(_05819_),
    .B2(_05057_),
    .X(_05820_));
 sky130_fd_sc_hd__mux2_2 _12641_ (.A0(\reg_gpout[2] ),
    .A1(clknet_1_1__leaf__05820_),
    .S(net45),
    .X(_05821_));
 sky130_fd_sc_hd__buf_1 _12642_ (.A(_05821_),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 _12643_ (.A(net22),
    .X(_05822_));
 sky130_fd_sc_hd__or2_1 _12644_ (.A(_05822_),
    .B(_05057_),
    .X(_05823_));
 sky130_fd_sc_hd__inv_2 _12645_ (.A(net25),
    .Y(_05824_));
 sky130_fd_sc_hd__nor2_1 _12646_ (.A(_05824_),
    .B(net26),
    .Y(_05825_));
 sky130_fd_sc_hd__nand2_1 _12647_ (.A(_05822_),
    .B(_05297_),
    .Y(_05826_));
 sky130_fd_sc_hd__mux4_1 _12648_ (.A0(_05382_),
    .A1(_05470_),
    .A2(_05551_),
    .A3(_05632_),
    .S0(_05822_),
    .S1(net25),
    .X(_05827_));
 sky130_fd_sc_hd__a32o_1 _12649_ (.A1(_05823_),
    .A2(_05825_),
    .A3(_05826_),
    .B1(_05827_),
    .B2(net26),
    .X(_05828_));
 sky130_fd_sc_hd__buf_2 _12650_ (.A(net24),
    .X(_05829_));
 sky130_fd_sc_hd__and4b_1 _12651_ (.A_N(net27),
    .B(_05828_),
    .C(net23),
    .D(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__a21o_1 _12652_ (.A1(net23),
    .A2(_05829_),
    .B1(net25),
    .X(_05831_));
 sky130_fd_sc_hd__nand2_1 _12653_ (.A(net26),
    .B(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hd__inv_2 _12654_ (.A(net23),
    .Y(_05833_));
 sky130_fd_sc_hd__mux4_1 _12655_ (.A0(_04687_),
    .A1(_05644_),
    .A2(_05645_),
    .A3(_04642_),
    .S0(_05822_),
    .S1(_05829_),
    .X(_05834_));
 sky130_fd_sc_hd__inv_2 _12656_ (.A(_05829_),
    .Y(_05835_));
 sky130_fd_sc_hd__mux4_1 _12657_ (.A0(_05650_),
    .A1(_05651_),
    .A2(_05652_),
    .A3(_05653_),
    .S0(_05822_),
    .S1(net25),
    .X(_05836_));
 sky130_fd_sc_hd__mux2_1 _12658_ (.A0(_05648_),
    .A1(_04657_),
    .S(_05822_),
    .X(_05837_));
 sky130_fd_sc_hd__or2_1 _12659_ (.A(_05829_),
    .B(_05837_),
    .X(_05838_));
 sky130_fd_sc_hd__o211a_1 _12660_ (.A1(_05835_),
    .A2(_05836_),
    .B1(_05838_),
    .C1(net23),
    .X(_05839_));
 sky130_fd_sc_hd__a21oi_1 _12661_ (.A1(_05833_),
    .A2(_05834_),
    .B1(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__nand2_1 _12662_ (.A(_05824_),
    .B(_05829_),
    .Y(_05841_));
 sky130_fd_sc_hd__nor2_1 _12663_ (.A(net23),
    .B(net22),
    .Y(_05842_));
 sky130_fd_sc_hd__and2_1 _12664_ (.A(_05833_),
    .B(net22),
    .X(_05843_));
 sky130_fd_sc_hd__a22oi_1 _12665_ (.A1(_05055_),
    .A2(_05842_),
    .B1(_05843_),
    .B2(net71),
    .Y(_05844_));
 sky130_fd_sc_hd__nor2_1 _12666_ (.A(_05833_),
    .B(_05822_),
    .Y(_05845_));
 sky130_fd_sc_hd__nor2_2 _12667_ (.A(net25),
    .B(net24),
    .Y(_05846_));
 sky130_fd_sc_hd__and2_1 _12668_ (.A(net23),
    .B(net22),
    .X(_05847_));
 sky130_fd_sc_hd__and3_1 _12669_ (.A(_05053_),
    .B(_05846_),
    .C(_05847_),
    .X(_05848_));
 sky130_fd_sc_hd__a22o_1 _12670_ (.A1(net41),
    .A2(_05845_),
    .B1(_05847_),
    .B2(_05263_),
    .X(_05849_));
 sky130_fd_sc_hd__a221o_1 _12671_ (.A1(net51),
    .A2(_05842_),
    .B1(_05843_),
    .B2(net40),
    .C1(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__nor2_1 _12672_ (.A(net27),
    .B(net26),
    .Y(_05851_));
 sky130_fd_sc_hd__a21o_1 _12673_ (.A1(_05711_),
    .A2(_05851_),
    .B1(net50),
    .X(_05852_));
 sky130_fd_sc_hd__a22o_1 _12674_ (.A1(net49),
    .A2(_05845_),
    .B1(_05847_),
    .B2(_05852_),
    .X(_05853_));
 sky130_fd_sc_hd__and2_1 _12675_ (.A(_05842_),
    .B(_05846_),
    .X(_05854_));
 sky130_fd_sc_hd__a32o_1 _12676_ (.A1(net46),
    .A2(_05843_),
    .A3(_05846_),
    .B1(_05854_),
    .B2(net43),
    .X(_05855_));
 sky130_fd_sc_hd__a31o_1 _12677_ (.A1(_05824_),
    .A2(_05829_),
    .A3(_05853_),
    .B1(_05855_),
    .X(_05856_));
 sky130_fd_sc_hd__a31o_1 _12678_ (.A1(net25),
    .A2(_05835_),
    .A3(_05850_),
    .B1(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__a311o_1 _12679_ (.A1(net44),
    .A2(_05845_),
    .A3(_05846_),
    .B1(_05848_),
    .C1(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__o21ba_1 _12680_ (.A1(_05841_),
    .A2(_05844_),
    .B1_N(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__o22ai_1 _12681_ (.A1(_05832_),
    .A2(_05840_),
    .B1(_05859_),
    .B2(net26),
    .Y(_05860_));
 sky130_fd_sc_hd__clkinv_2 _12682_ (.A(_05711_),
    .Y(_05861_));
 sky130_fd_sc_hd__and4bb_1 _12683_ (.A_N(_05861_),
    .B_N(_05841_),
    .C(_05847_),
    .D(_05851_),
    .X(_05862_));
 sky130_fd_sc_hd__a21o_1 _12684_ (.A1(net25),
    .A2(_05829_),
    .B1(net26),
    .X(_05863_));
 sky130_fd_sc_hd__and3_1 _12685_ (.A(net27),
    .B(_05832_),
    .C(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__mux4_1 _12686_ (.A0(_04589_),
    .A1(_04704_),
    .A2(_04419_),
    .A3(_03973_),
    .S0(_05822_),
    .S1(net23),
    .X(_05865_));
 sky130_fd_sc_hd__mux4_1 _12687_ (.A0(_03969_),
    .A1(_04575_),
    .A2(_04452_),
    .A3(_04628_),
    .S0(_05822_),
    .S1(net23),
    .X(_05866_));
 sky130_fd_sc_hd__mux2_1 _12688_ (.A0(_03975_),
    .A1(_04420_),
    .S(_05822_),
    .X(_05867_));
 sky130_fd_sc_hd__mux2_1 _12689_ (.A0(_05866_),
    .A1(_05867_),
    .S(_05824_),
    .X(_05868_));
 sky130_fd_sc_hd__mux2_1 _12690_ (.A0(_05865_),
    .A1(_05868_),
    .S(_05829_),
    .X(_05869_));
 sky130_fd_sc_hd__a22o_1 _12691_ (.A1(net53),
    .A2(_05843_),
    .B1(_05845_),
    .B2(net55),
    .X(_05870_));
 sky130_fd_sc_hd__a21o_1 _12692_ (.A1(net52),
    .A2(_05842_),
    .B1(_05870_),
    .X(_05871_));
 sky130_fd_sc_hd__a31o_1 _12693_ (.A1(net48),
    .A2(_05833_),
    .A3(_05846_),
    .B1(_05854_),
    .X(_05872_));
 sky130_fd_sc_hd__a31o_1 _12694_ (.A1(\gpout3.clk_div[1] ),
    .A2(_05846_),
    .A3(_05847_),
    .B1(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__a31o_2 _12695_ (.A1(clknet_1_0__leaf__04634_),
    .A2(_05845_),
    .A3(_05846_),
    .B1(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__a31o_2 _12696_ (.A1(_05824_),
    .A2(_05829_),
    .A3(_05871_),
    .B1(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__a22o_2 _12697_ (.A1(_05864_),
    .A2(_05869_),
    .B1(_05875_),
    .B2(_05851_),
    .X(_05876_));
 sky130_fd_sc_hd__a211o_2 _12698_ (.A1(net27),
    .A2(_05860_),
    .B1(_05862_),
    .C1(_05876_),
    .X(_05877_));
 sky130_fd_sc_hd__nand2_1 _12699_ (.A(_05851_),
    .B(_05854_),
    .Y(_05878_));
 sky130_fd_sc_hd__o22a_2 _12700_ (.A1(_05830_),
    .A2(_05877_),
    .B1(_05878_),
    .B2(_05298_),
    .X(_05879_));
 sky130_fd_sc_hd__mux2_2 _12701_ (.A0(\reg_gpout[3] ),
    .A1(clknet_1_0__leaf__05879_),
    .S(net45),
    .X(_05880_));
 sky130_fd_sc_hd__buf_1 _12702_ (.A(_05880_),
    .X(net59));
 sky130_fd_sc_hd__buf_2 _12703_ (.A(net28),
    .X(_05881_));
 sky130_fd_sc_hd__or2_1 _12704_ (.A(_05881_),
    .B(_05057_),
    .X(_05882_));
 sky130_fd_sc_hd__nand2_1 _12705_ (.A(_05881_),
    .B(_05297_),
    .Y(_05883_));
 sky130_fd_sc_hd__inv_2 _12706_ (.A(net31),
    .Y(_05884_));
 sky130_fd_sc_hd__nor2_1 _12707_ (.A(_05884_),
    .B(net32),
    .Y(_05885_));
 sky130_fd_sc_hd__mux4_1 _12708_ (.A0(_05382_),
    .A1(_05470_),
    .A2(_05551_),
    .A3(_05632_),
    .S0(_05881_),
    .S1(net31),
    .X(_05886_));
 sky130_fd_sc_hd__a32o_1 _12709_ (.A1(_05882_),
    .A2(_05883_),
    .A3(_05885_),
    .B1(_05886_),
    .B2(net32),
    .X(_05887_));
 sky130_fd_sc_hd__buf_2 _12710_ (.A(net29),
    .X(_05888_));
 sky130_fd_sc_hd__buf_2 _12711_ (.A(net30),
    .X(_05889_));
 sky130_fd_sc_hd__and4b_1 _12712_ (.A_N(net33),
    .B(_05887_),
    .C(_05888_),
    .D(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__a21oi_1 _12713_ (.A1(_05888_),
    .A2(_05889_),
    .B1(net31),
    .Y(_05891_));
 sky130_fd_sc_hd__a22o_1 _12714_ (.A1(_05889_),
    .A2(_05885_),
    .B1(_05891_),
    .B2(net32),
    .X(_05892_));
 sky130_fd_sc_hd__mux4_1 _12715_ (.A0(_04589_),
    .A1(_04704_),
    .A2(_04419_),
    .A3(_03973_),
    .S0(_05881_),
    .S1(_05888_),
    .X(_05893_));
 sky130_fd_sc_hd__mux4_1 _12716_ (.A0(_03969_),
    .A1(_04575_),
    .A2(_04452_),
    .A3(_04628_),
    .S0(net28),
    .S1(net29),
    .X(_05894_));
 sky130_fd_sc_hd__mux2_1 _12717_ (.A0(_03975_),
    .A1(_04420_),
    .S(net28),
    .X(_05895_));
 sky130_fd_sc_hd__mux2_1 _12718_ (.A0(_05894_),
    .A1(_05895_),
    .S(_05884_),
    .X(_05896_));
 sky130_fd_sc_hd__mux2_1 _12719_ (.A0(_05893_),
    .A1(_05896_),
    .S(_05889_),
    .X(_05897_));
 sky130_fd_sc_hd__and3_1 _12720_ (.A(net33),
    .B(_05892_),
    .C(_05897_),
    .X(_05898_));
 sky130_fd_sc_hd__inv_2 _12721_ (.A(net29),
    .Y(_05899_));
 sky130_fd_sc_hd__mux4_1 _12722_ (.A0(_04687_),
    .A1(_04653_),
    .A2(_05645_),
    .A3(_04642_),
    .S0(_05881_),
    .S1(_05889_),
    .X(_05900_));
 sky130_fd_sc_hd__inv_2 _12723_ (.A(_05889_),
    .Y(_05901_));
 sky130_fd_sc_hd__mux4_1 _12724_ (.A0(\gpout0.vpos[0] ),
    .A1(_05651_),
    .A2(_05652_),
    .A3(_05653_),
    .S0(net28),
    .S1(net31),
    .X(_05902_));
 sky130_fd_sc_hd__or2_1 _12725_ (.A(_05901_),
    .B(_05902_),
    .X(_05903_));
 sky130_fd_sc_hd__mux2_1 _12726_ (.A0(_05648_),
    .A1(_04657_),
    .S(net28),
    .X(_05904_));
 sky130_fd_sc_hd__o21a_1 _12727_ (.A1(_05889_),
    .A2(_05904_),
    .B1(_05888_),
    .X(_05905_));
 sky130_fd_sc_hd__a22o_1 _12728_ (.A1(_05899_),
    .A2(_05900_),
    .B1(_05903_),
    .B2(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__and4b_1 _12729_ (.A_N(_05891_),
    .B(_05906_),
    .C(net32),
    .D(net33),
    .X(_05907_));
 sky130_fd_sc_hd__mux4_1 _12730_ (.A0(net51),
    .A1(net41),
    .A2(net40),
    .A3(_05263_),
    .S0(_05888_),
    .S1(_05881_),
    .X(_05908_));
 sky130_fd_sc_hd__nor2_2 _12731_ (.A(net31),
    .B(net30),
    .Y(_05909_));
 sky130_fd_sc_hd__nor2_1 _12732_ (.A(_05899_),
    .B(_05881_),
    .Y(_05910_));
 sky130_fd_sc_hd__nor2_1 _12733_ (.A(net32),
    .B(net33),
    .Y(_05911_));
 sky130_fd_sc_hd__a21o_1 _12734_ (.A1(_05711_),
    .A2(_05911_),
    .B1(net50),
    .X(_05912_));
 sky130_fd_sc_hd__and3_1 _12735_ (.A(_05888_),
    .B(net28),
    .C(_05912_),
    .X(_05913_));
 sky130_fd_sc_hd__a21oi_1 _12736_ (.A1(net49),
    .A2(_05910_),
    .B1(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__nor2_1 _12737_ (.A(net31),
    .B(_05914_),
    .Y(_05915_));
 sky130_fd_sc_hd__a211o_1 _12738_ (.A1(_05901_),
    .A2(_05908_),
    .B1(_05909_),
    .C1(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__and4_1 _12739_ (.A(_05888_),
    .B(_05881_),
    .C(_05884_),
    .D(_05889_),
    .X(_05917_));
 sky130_fd_sc_hd__and2b_1 _12740_ (.A_N(net32),
    .B(net33),
    .X(_05918_));
 sky130_fd_sc_hd__a31o_1 _12741_ (.A1(_05711_),
    .A2(_05911_),
    .A3(_05917_),
    .B1(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__and2_1 _12742_ (.A(_05899_),
    .B(net28),
    .X(_05920_));
 sky130_fd_sc_hd__nor2_1 _12743_ (.A(net29),
    .B(net28),
    .Y(_05921_));
 sky130_fd_sc_hd__or2_1 _12744_ (.A(net31),
    .B(net30),
    .X(_05922_));
 sky130_fd_sc_hd__a221o_1 _12745_ (.A1(net46),
    .A2(_05920_),
    .B1(_05921_),
    .B2(net43),
    .C1(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__and2_1 _12746_ (.A(net52),
    .B(_05921_),
    .X(_05924_));
 sky130_fd_sc_hd__a221o_1 _12747_ (.A1(net55),
    .A2(_05910_),
    .B1(_05920_),
    .B2(net53),
    .C1(_05924_),
    .X(_05925_));
 sky130_fd_sc_hd__a211oi_1 _12748_ (.A1(_04643_),
    .A2(net28),
    .B1(_05922_),
    .C1(_05888_),
    .Y(_05926_));
 sky130_fd_sc_hd__a41o_1 _12749_ (.A1(_05888_),
    .A2(_05881_),
    .A3(\gpout4.clk_div[1] ),
    .A4(_05909_),
    .B1(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__a31o_2 _12750_ (.A1(clknet_1_0__leaf__04634_),
    .A2(_05910_),
    .A3(_05909_),
    .B1(_05927_),
    .X(_05928_));
 sky130_fd_sc_hd__a31o_2 _12751_ (.A1(_05884_),
    .A2(_05889_),
    .A3(_05925_),
    .B1(_05928_),
    .X(_05929_));
 sky130_fd_sc_hd__a32o_2 _12752_ (.A1(_05916_),
    .A2(_05919_),
    .A3(_05923_),
    .B1(_05929_),
    .B2(_05911_),
    .X(_05930_));
 sky130_fd_sc_hd__a22o_1 _12753_ (.A1(net71),
    .A2(_05920_),
    .B1(_05921_),
    .B2(_05055_),
    .X(_05931_));
 sky130_fd_sc_hd__and3_1 _12754_ (.A(_05884_),
    .B(_05889_),
    .C(_05931_),
    .X(_05932_));
 sky130_fd_sc_hd__and4_1 _12755_ (.A(_05888_),
    .B(_05881_),
    .C(_05053_),
    .D(_05909_),
    .X(_05933_));
 sky130_fd_sc_hd__a31o_1 _12756_ (.A1(net44),
    .A2(_05910_),
    .A3(_05909_),
    .B1(_05933_),
    .X(_05934_));
 sky130_fd_sc_hd__o21a_1 _12757_ (.A1(_05932_),
    .A2(_05934_),
    .B1(_05918_),
    .X(_05935_));
 sky130_fd_sc_hd__or4_2 _12758_ (.A(_05898_),
    .B(_05907_),
    .C(_05930_),
    .D(_05935_),
    .X(_05936_));
 sky130_fd_sc_hd__nand3_1 _12759_ (.A(_05911_),
    .B(_05921_),
    .C(_05909_),
    .Y(_05937_));
 sky130_fd_sc_hd__o22a_2 _12760_ (.A1(_05890_),
    .A2(_05936_),
    .B1(_05937_),
    .B2(_05551_),
    .X(_05938_));
 sky130_fd_sc_hd__mux2_2 _12761_ (.A0(\reg_gpout[4] ),
    .A1(clknet_1_1__leaf__05938_),
    .S(net45),
    .X(_05939_));
 sky130_fd_sc_hd__buf_1 _12762_ (.A(_05939_),
    .X(net60));
 sky130_fd_sc_hd__or2_1 _12763_ (.A(net37),
    .B(net36),
    .X(_05940_));
 sky130_fd_sc_hd__nor2_2 _12764_ (.A(net35),
    .B(net34),
    .Y(_05941_));
 sky130_fd_sc_hd__nor2_1 _12765_ (.A(net38),
    .B(net39),
    .Y(_05942_));
 sky130_fd_sc_hd__nand2_1 _12766_ (.A(_05941_),
    .B(_05942_),
    .Y(_05943_));
 sky130_fd_sc_hd__and2b_1 _12767_ (.A_N(net35),
    .B(net34),
    .X(_05944_));
 sky130_fd_sc_hd__and2b_1 _12768_ (.A_N(net34),
    .B(net35),
    .X(_05945_));
 sky130_fd_sc_hd__buf_2 _12769_ (.A(net35),
    .X(_05946_));
 sky130_fd_sc_hd__and3_1 _12770_ (.A(net50),
    .B(_05946_),
    .C(net34),
    .X(_05947_));
 sky130_fd_sc_hd__buf_2 _12771_ (.A(net36),
    .X(_05948_));
 sky130_fd_sc_hd__inv_2 _12772_ (.A(_05948_),
    .Y(_05949_));
 sky130_fd_sc_hd__a211o_1 _12773_ (.A1(net49),
    .A2(_05945_),
    .B1(_05947_),
    .C1(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__a221o_1 _12774_ (.A1(net71),
    .A2(_05944_),
    .B1(_05941_),
    .B2(_05055_),
    .C1(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__inv_2 _12775_ (.A(net37),
    .Y(_05952_));
 sky130_fd_sc_hd__and3_1 _12776_ (.A(_05946_),
    .B(net34),
    .C(_05053_),
    .X(_05953_));
 sky130_fd_sc_hd__a221o_1 _12777_ (.A1(net44),
    .A2(_05945_),
    .B1(_05941_),
    .B2(net43),
    .C1(_05940_),
    .X(_05954_));
 sky130_fd_sc_hd__a211o_1 _12778_ (.A1(net46),
    .A2(_05944_),
    .B1(_05953_),
    .C1(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__a221o_1 _12779_ (.A1(net40),
    .A2(_05944_),
    .B1(_05941_),
    .B2(net51),
    .C1(_05952_),
    .X(_05956_));
 sky130_fd_sc_hd__o211a_1 _12780_ (.A1(_05952_),
    .A2(_05949_),
    .B1(_05955_),
    .C1(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__clkbuf_4 _12781_ (.A(net34),
    .X(_05958_));
 sky130_fd_sc_hd__mux4_1 _12782_ (.A0(_03969_),
    .A1(_04575_),
    .A2(_04452_),
    .A3(_04628_),
    .S0(_05958_),
    .S1(_05946_),
    .X(_05959_));
 sky130_fd_sc_hd__a31o_1 _12783_ (.A1(net37),
    .A2(_05948_),
    .A3(_05959_),
    .B1(net38),
    .X(_05960_));
 sky130_fd_sc_hd__a21o_1 _12784_ (.A1(_05951_),
    .A2(_05957_),
    .B1(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__mux2_1 _12785_ (.A0(_05650_),
    .A1(_05651_),
    .S(_05958_),
    .X(_05962_));
 sky130_fd_sc_hd__mux4_1 _12786_ (.A0(_04589_),
    .A1(_04704_),
    .A2(_04419_),
    .A3(_03973_),
    .S0(net34),
    .S1(net35),
    .X(_05963_));
 sky130_fd_sc_hd__a22o_1 _12787_ (.A1(_04420_),
    .A2(_05944_),
    .B1(_05941_),
    .B2(_03975_),
    .X(_05964_));
 sky130_fd_sc_hd__mux2_1 _12788_ (.A0(_05963_),
    .A1(_05964_),
    .S(_05948_),
    .X(_05965_));
 sky130_fd_sc_hd__a31o_1 _12789_ (.A1(_05946_),
    .A2(_05948_),
    .A3(_05962_),
    .B1(_05965_),
    .X(_05966_));
 sky130_fd_sc_hd__mux2_1 _12790_ (.A0(_05652_),
    .A1(_05653_),
    .S(net34),
    .X(_05967_));
 sky130_fd_sc_hd__nand2_1 _12791_ (.A(_05948_),
    .B(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__nor2_1 _12792_ (.A(_05648_),
    .B(_05958_),
    .Y(_05969_));
 sky130_fd_sc_hd__a211o_1 _12793_ (.A1(_04731_),
    .A2(_05958_),
    .B1(_05948_),
    .C1(_05969_),
    .X(_05970_));
 sky130_fd_sc_hd__mux4_1 _12794_ (.A0(_04687_),
    .A1(_04653_),
    .A2(_05645_),
    .A3(_04642_),
    .S0(net34),
    .S1(_05948_),
    .X(_05971_));
 sky130_fd_sc_hd__o21ai_1 _12795_ (.A1(_05946_),
    .A2(_05971_),
    .B1(net37),
    .Y(_05972_));
 sky130_fd_sc_hd__a31o_1 _12796_ (.A1(_05946_),
    .A2(_05968_),
    .A3(_05970_),
    .B1(_05972_),
    .X(_05973_));
 sky130_fd_sc_hd__nand2_1 _12797_ (.A(net38),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__a21o_1 _12798_ (.A1(_05952_),
    .A2(_05966_),
    .B1(_05974_),
    .X(_05975_));
 sky130_fd_sc_hd__or2_1 _12799_ (.A(_05958_),
    .B(_05057_),
    .X(_05976_));
 sky130_fd_sc_hd__nor2_1 _12800_ (.A(_05952_),
    .B(net38),
    .Y(_05977_));
 sky130_fd_sc_hd__nand2_1 _12801_ (.A(_05958_),
    .B(_05297_),
    .Y(_05978_));
 sky130_fd_sc_hd__mux4_1 _12802_ (.A0(_05382_),
    .A1(_05470_),
    .A2(_05551_),
    .A3(_05632_),
    .S0(_05958_),
    .S1(net37),
    .X(_05979_));
 sky130_fd_sc_hd__a32o_1 _12803_ (.A1(_05976_),
    .A2(_05977_),
    .A3(_05978_),
    .B1(_05979_),
    .B2(net38),
    .X(_05980_));
 sky130_fd_sc_hd__and4b_1 _12804_ (.A_N(net39),
    .B(_05980_),
    .C(_05946_),
    .D(_05948_),
    .X(_05981_));
 sky130_fd_sc_hd__a22o_1 _12805_ (.A1(net55),
    .A2(_05945_),
    .B1(_05941_),
    .B2(net52),
    .X(_05982_));
 sky130_fd_sc_hd__a21o_1 _12806_ (.A1(net53),
    .A2(_05944_),
    .B1(_05982_),
    .X(_05983_));
 sky130_fd_sc_hd__and3_1 _12807_ (.A(_05711_),
    .B(_05952_),
    .C(_05948_),
    .X(_05984_));
 sky130_fd_sc_hd__a31o_1 _12808_ (.A1(_05952_),
    .A2(_05949_),
    .A3(\gpout5.clk_div[1] ),
    .B1(_05984_),
    .X(_05985_));
 sky130_fd_sc_hd__a211oi_2 _12809_ (.A1(net126),
    .A2(_05946_),
    .B1(_05958_),
    .C1(_05940_),
    .Y(_05986_));
 sky130_fd_sc_hd__a31o_2 _12810_ (.A1(_05946_),
    .A2(_05958_),
    .A3(_05985_),
    .B1(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__a31o_2 _12811_ (.A1(_05952_),
    .A2(_05948_),
    .A3(_05983_),
    .B1(_05987_),
    .X(_05988_));
 sky130_fd_sc_hd__mux2_1 _12812_ (.A0(net41),
    .A1(_05263_),
    .S(_05958_),
    .X(_05989_));
 sky130_fd_sc_hd__and4_1 _12813_ (.A(_05949_),
    .B(net39),
    .C(_05977_),
    .D(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__a22o_2 _12814_ (.A1(_05988_),
    .A2(_05942_),
    .B1(_05990_),
    .B2(_05946_),
    .X(_05991_));
 sky130_fd_sc_hd__a311o_2 _12815_ (.A1(net39),
    .A2(_05961_),
    .A3(_05975_),
    .B1(_05981_),
    .C1(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__o31a_2 _12816_ (.A1(_05632_),
    .A2(_05940_),
    .A3(_05943_),
    .B1(_05992_),
    .X(_05993_));
 sky130_fd_sc_hd__mux2_2 _12817_ (.A0(\reg_gpout[5] ),
    .A1(clknet_1_0__leaf__05993_),
    .S(net45),
    .X(_05994_));
 sky130_fd_sc_hd__buf_1 _12818_ (.A(_05994_),
    .X(net61));
 sky130_fd_sc_hd__and2_1 _12819_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(_05995_));
 sky130_fd_sc_hd__nand2_1 _12820_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_05996_));
 sky130_fd_sc_hd__or2_1 _12821_ (.A(\rbzero.debug_overlay.facingY[0] ),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .X(_05997_));
 sky130_fd_sc_hd__nand3_1 _12822_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .C(_05997_),
    .Y(_05998_));
 sky130_fd_sc_hd__xnor2_1 _12823_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_05999_));
 sky130_fd_sc_hd__and2_1 _12824_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_06000_));
 sky130_fd_sc_hd__nor2_1 _12825_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_06001_));
 sky130_fd_sc_hd__or3_1 _12826_ (.A(_05999_),
    .B(_06000_),
    .C(_06001_),
    .X(_06002_));
 sky130_fd_sc_hd__nand2_1 _12827_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_06003_));
 sky130_fd_sc_hd__or2_1 _12828_ (.A(\rbzero.debug_overlay.facingY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_06004_));
 sky130_fd_sc_hd__and2_1 _12829_ (.A(_06003_),
    .B(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__nor2_1 _12830_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_06006_));
 sky130_fd_sc_hd__and2_1 _12831_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_06007_));
 sky130_fd_sc_hd__nor2_1 _12832_ (.A(_06006_),
    .B(_06007_),
    .Y(_06008_));
 sky130_fd_sc_hd__nand2_1 _12833_ (.A(_06005_),
    .B(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__or2_1 _12834_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .X(_06010_));
 sky130_fd_sc_hd__and2_1 _12835_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_06011_));
 sky130_fd_sc_hd__nor2_1 _12836_ (.A(\rbzero.debug_overlay.facingY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_06012_));
 sky130_fd_sc_hd__nor2_1 _12837_ (.A(_06011_),
    .B(_06012_),
    .Y(_06013_));
 sky130_fd_sc_hd__xor2_2 _12838_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_06014_));
 sky130_fd_sc_hd__and2_1 _12839_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_06015_));
 sky130_fd_sc_hd__a31o_1 _12840_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A3(_06014_),
    .B1(_06015_),
    .X(_06016_));
 sky130_fd_sc_hd__a221o_1 _12841_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1(_06013_),
    .B2(_06016_),
    .C1(_06011_),
    .X(_06017_));
 sky130_fd_sc_hd__or4bb_1 _12842_ (.A(_06002_),
    .B(_06009_),
    .C_N(_06010_),
    .D_N(_06017_),
    .X(_06018_));
 sky130_fd_sc_hd__nor2_1 _12843_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_06019_));
 sky130_fd_sc_hd__nand2_1 _12844_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_06020_));
 sky130_fd_sc_hd__nand2_1 _12845_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .Y(_06021_));
 sky130_fd_sc_hd__a211o_1 _12846_ (.A1(_06003_),
    .A2(_06021_),
    .B1(_06006_),
    .C1(_06002_),
    .X(_06022_));
 sky130_fd_sc_hd__nand2_1 _12847_ (.A(\rbzero.debug_overlay.facingY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_06023_));
 sky130_fd_sc_hd__o211a_1 _12848_ (.A1(_06019_),
    .A2(_06020_),
    .B1(_06022_),
    .C1(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__nand2_1 _12849_ (.A(_05997_),
    .B(_05996_),
    .Y(_06025_));
 sky130_fd_sc_hd__nand2_1 _12850_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_06026_));
 sky130_fd_sc_hd__or2_1 _12851_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_06027_));
 sky130_fd_sc_hd__nand2_1 _12852_ (.A(_06026_),
    .B(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__a211o_1 _12853_ (.A1(_06018_),
    .A2(_06024_),
    .B1(_06025_),
    .C1(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__nand2_1 _12854_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_06030_));
 sky130_fd_sc_hd__nor2_1 _12855_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_06031_));
 sky130_fd_sc_hd__a41o_2 _12856_ (.A1(_05996_),
    .A2(_05998_),
    .A3(_06029_),
    .A4(_06030_),
    .B1(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__or2_2 _12857_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .X(_06033_));
 sky130_fd_sc_hd__o21ai_4 _12858_ (.A1(_05995_),
    .A2(_06032_),
    .B1(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__nand2_1 _12859_ (.A(\rbzero.debug_overlay.facingY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_06035_));
 sky130_fd_sc_hd__nand2_1 _12860_ (.A(_06033_),
    .B(_06035_),
    .Y(_06036_));
 sky130_fd_sc_hd__xor2_2 _12861_ (.A(_06032_),
    .B(_06036_),
    .X(_06037_));
 sky130_fd_sc_hd__and2b_1 _12862_ (.A_N(_06031_),
    .B(_06030_),
    .X(_06038_));
 sky130_fd_sc_hd__a31oi_2 _12863_ (.A1(_05996_),
    .A2(_05998_),
    .A3(_06029_),
    .B1(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__and4_1 _12864_ (.A(_05996_),
    .B(_05998_),
    .C(_06029_),
    .D(_06038_),
    .X(_06040_));
 sky130_fd_sc_hd__or2_1 _12865_ (.A(_06039_),
    .B(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__inv_2 _12866_ (.A(_06026_),
    .Y(_06042_));
 sky130_fd_sc_hd__a21oi_2 _12867_ (.A1(_06018_),
    .A2(_06024_),
    .B1(_06028_),
    .Y(_06043_));
 sky130_fd_sc_hd__o21bai_2 _12868_ (.A1(_06042_),
    .A2(_06043_),
    .B1_N(_06025_),
    .Y(_06044_));
 sky130_fd_sc_hd__or3b_1 _12869_ (.A(_06042_),
    .B(_06043_),
    .C_N(_06025_),
    .X(_06045_));
 sky130_fd_sc_hd__nand3_1 _12870_ (.A(_06010_),
    .B(_06017_),
    .C(_06005_),
    .Y(_06046_));
 sky130_fd_sc_hd__or2_1 _12871_ (.A(_06000_),
    .B(_06001_),
    .X(_06047_));
 sky130_fd_sc_hd__a311o_1 _12872_ (.A1(_06003_),
    .A2(_06046_),
    .A3(_06021_),
    .B1(_06006_),
    .C1(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__or2_1 _12873_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_06049_));
 sky130_fd_sc_hd__a32o_1 _12874_ (.A1(_06010_),
    .A2(_06017_),
    .A3(_06005_),
    .B1(\rbzero.wall_tracer.rayAddendY[3] ),
    .B2(\rbzero.debug_overlay.facingY[-5] ),
    .X(_06050_));
 sky130_fd_sc_hd__nor2_1 _12875_ (.A(_06000_),
    .B(_06001_),
    .Y(_06051_));
 sky130_fd_sc_hd__a211o_1 _12876_ (.A1(_06049_),
    .A2(_06050_),
    .B1(_06007_),
    .C1(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__and2_1 _12877_ (.A(_06048_),
    .B(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__and3_1 _12878_ (.A(_06028_),
    .B(_06018_),
    .C(_06024_),
    .X(_06054_));
 sky130_fd_sc_hd__nor2_1 _12879_ (.A(_06043_),
    .B(_06054_),
    .Y(_06055_));
 sky130_fd_sc_hd__xor2_1 _12880_ (.A(_06008_),
    .B(_06050_),
    .X(_06056_));
 sky130_fd_sc_hd__a21o_1 _12881_ (.A1(_06010_),
    .A2(_06017_),
    .B1(_06005_),
    .X(_06057_));
 sky130_fd_sc_hd__and2_1 _12882_ (.A(_06046_),
    .B(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__nand2_1 _12883_ (.A(\rbzero.debug_overlay.facingY[-6] ),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_06059_));
 sky130_fd_sc_hd__nand2_1 _12884_ (.A(_06010_),
    .B(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__a21o_1 _12885_ (.A1(_06013_),
    .A2(_06016_),
    .B1(_06011_),
    .X(_06061_));
 sky130_fd_sc_hd__xnor2_1 _12886_ (.A(_06060_),
    .B(_06061_),
    .Y(_06062_));
 sky130_fd_sc_hd__xor2_2 _12887_ (.A(_06013_),
    .B(_06016_),
    .X(_06063_));
 sky130_fd_sc_hd__nand2_1 _12888_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_06064_));
 sky130_fd_sc_hd__xnor2_2 _12889_ (.A(_06064_),
    .B(_06014_),
    .Y(_06065_));
 sky130_fd_sc_hd__xor2_2 _12890_ (.A(\rbzero.debug_overlay.facingY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_06066_));
 sky130_fd_sc_hd__or4_1 _12891_ (.A(\rbzero.wall_tracer.rayAddendY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .C(_06065_),
    .D(_06066_),
    .X(_06067_));
 sky130_fd_sc_hd__or4_1 _12892_ (.A(_06058_),
    .B(_06062_),
    .C(_06063_),
    .D(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__or3_1 _12893_ (.A(_06055_),
    .B(_06056_),
    .C(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__a211o_1 _12894_ (.A1(_06044_),
    .A2(_06045_),
    .B1(_06053_),
    .C1(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__a21o_1 _12895_ (.A1(_06020_),
    .A2(_06048_),
    .B1(_05999_),
    .X(_06071_));
 sky130_fd_sc_hd__nand3_1 _12896_ (.A(_05999_),
    .B(_06020_),
    .C(_06048_),
    .Y(_06072_));
 sky130_fd_sc_hd__nand2_1 _12897_ (.A(_06071_),
    .B(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__or4b_2 _12898_ (.A(_06037_),
    .B(_06041_),
    .C(_06070_),
    .D_N(_06073_),
    .X(_06074_));
 sky130_fd_sc_hd__nand2_1 _12899_ (.A(_06034_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__buf_4 _12900_ (.A(_06075_),
    .X(_06076_));
 sky130_fd_sc_hd__clkbuf_4 _12901_ (.A(_06076_),
    .X(_06077_));
 sky130_fd_sc_hd__buf_2 _12902_ (.A(_06077_),
    .X(_06078_));
 sky130_fd_sc_hd__o21a_1 _12903_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(\rbzero.wall_tracer.mapY[5] ),
    .B1(_06078_),
    .X(_06079_));
 sky130_fd_sc_hd__inv_2 _12904_ (.A(\rbzero.wall_tracer.mapY[5] ),
    .Y(_06080_));
 sky130_fd_sc_hd__xnor2_1 _12905_ (.A(_06080_),
    .B(_06077_),
    .Y(_06081_));
 sky130_fd_sc_hd__nand2_1 _12906_ (.A(\rbzero.map_rom.i_row[4] ),
    .B(_06077_),
    .Y(_06082_));
 sky130_fd_sc_hd__or2_1 _12907_ (.A(\rbzero.map_rom.i_row[4] ),
    .B(_06077_),
    .X(_06083_));
 sky130_fd_sc_hd__nand2_1 _12908_ (.A(\rbzero.map_rom.a6 ),
    .B(_06077_),
    .Y(_06084_));
 sky130_fd_sc_hd__inv_2 _12909_ (.A(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__inv_2 _12910_ (.A(\rbzero.map_rom.b6 ),
    .Y(_06086_));
 sky130_fd_sc_hd__inv_2 _12911_ (.A(_06076_),
    .Y(_06087_));
 sky130_fd_sc_hd__buf_2 _12912_ (.A(\rbzero.map_rom.d6 ),
    .X(_06088_));
 sky130_fd_sc_hd__clkinv_2 _12913_ (.A(\rbzero.map_rom.c6 ),
    .Y(_06089_));
 sky130_fd_sc_hd__xnor2_1 _12914_ (.A(_06089_),
    .B(_06076_),
    .Y(_06090_));
 sky130_fd_sc_hd__and2_1 _12915_ (.A(_06088_),
    .B(_06090_),
    .X(_06091_));
 sky130_fd_sc_hd__a21o_1 _12916_ (.A1(\rbzero.map_rom.c6 ),
    .A2(_06077_),
    .B1(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__xnor2_1 _12917_ (.A(_06086_),
    .B(_06076_),
    .Y(_06093_));
 sky130_fd_sc_hd__nand2_1 _12918_ (.A(_06092_),
    .B(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__o21ai_1 _12919_ (.A1(_06086_),
    .A2(_06087_),
    .B1(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__or2_1 _12920_ (.A(\rbzero.map_rom.a6 ),
    .B(_06077_),
    .X(_06096_));
 sky130_fd_sc_hd__o21a_1 _12921_ (.A1(_06085_),
    .A2(_06095_),
    .B1(_06096_),
    .X(_06097_));
 sky130_fd_sc_hd__and3_1 _12922_ (.A(_06082_),
    .B(_06083_),
    .C(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__and2_1 _12923_ (.A(_06081_),
    .B(_06098_),
    .X(_06099_));
 sky130_fd_sc_hd__xor2_1 _12924_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(_06077_),
    .X(_06100_));
 sky130_fd_sc_hd__o21ai_1 _12925_ (.A1(_06079_),
    .A2(_06099_),
    .B1(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__or3_1 _12926_ (.A(_06100_),
    .B(_06079_),
    .C(_06099_),
    .X(_06102_));
 sky130_fd_sc_hd__or3b_2 _12927_ (.A(_04429_),
    .B(_04430_),
    .C_N(\rbzero.trace_state[3] ),
    .X(_06103_));
 sky130_fd_sc_hd__buf_4 _12928_ (.A(_06103_),
    .X(_06104_));
 sky130_fd_sc_hd__buf_6 _12929_ (.A(_06104_),
    .X(_06105_));
 sky130_fd_sc_hd__nor3b_2 _12930_ (.A(_04429_),
    .B(_04430_),
    .C_N(\rbzero.trace_state[3] ),
    .Y(_06106_));
 sky130_fd_sc_hd__inv_2 _12931_ (.A(\rbzero.map_rom.a6 ),
    .Y(_06107_));
 sky130_fd_sc_hd__inv_2 _12932_ (.A(\rbzero.map_rom.f4 ),
    .Y(_06108_));
 sky130_fd_sc_hd__a22o_1 _12933_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_06108_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_04673_),
    .X(_06109_));
 sky130_fd_sc_hd__a221o_1 _12934_ (.A1(_04679_),
    .A2(\rbzero.map_rom.f4 ),
    .B1(_06107_),
    .B2(\rbzero.debug_overlay.playerY[3] ),
    .C1(_06109_),
    .X(_06110_));
 sky130_fd_sc_hd__inv_2 _12935_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .Y(_06111_));
 sky130_fd_sc_hd__inv_2 _12936_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .Y(_06112_));
 sky130_fd_sc_hd__clkbuf_4 _12937_ (.A(\rbzero.map_rom.f3 ),
    .X(_06113_));
 sky130_fd_sc_hd__inv_2 _12938_ (.A(\rbzero.debug_overlay.playerY[5] ),
    .Y(_06114_));
 sky130_fd_sc_hd__a22o_1 _12939_ (.A1(_04671_),
    .A2(_06113_),
    .B1(\rbzero.wall_tracer.mapY[5] ),
    .B2(_06114_),
    .X(_06115_));
 sky130_fd_sc_hd__a221o_1 _12940_ (.A1(_06111_),
    .A2(\rbzero.map_rom.c6 ),
    .B1(\rbzero.map_rom.b6 ),
    .B2(_06112_),
    .C1(_06115_),
    .X(_06116_));
 sky130_fd_sc_hd__clkinv_2 _12941_ (.A(\rbzero.map_rom.f3 ),
    .Y(_06117_));
 sky130_fd_sc_hd__nor2_1 _12942_ (.A(_06111_),
    .B(\rbzero.map_rom.c6 ),
    .Y(_06118_));
 sky130_fd_sc_hd__a221o_1 _12943_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_06117_),
    .B1(_06080_),
    .B2(\rbzero.debug_overlay.playerY[5] ),
    .C1(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__clkinv_2 _12944_ (.A(\rbzero.map_rom.f2 ),
    .Y(_06120_));
 sky130_fd_sc_hd__inv_2 _12945_ (.A(\rbzero.map_rom.i_row[4] ),
    .Y(_06121_));
 sky130_fd_sc_hd__xor2_1 _12946_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(\rbzero.map_rom.f1 ),
    .X(_06122_));
 sky130_fd_sc_hd__a221o_1 _12947_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_06120_),
    .B1(_06121_),
    .B2(\rbzero.debug_overlay.playerY[4] ),
    .C1(_06122_),
    .X(_06123_));
 sky130_fd_sc_hd__or4_1 _12948_ (.A(_06110_),
    .B(_06116_),
    .C(_06119_),
    .D(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__or4_1 _12949_ (.A(\rbzero.wall_tracer.mapY[6] ),
    .B(\rbzero.wall_tracer.mapY[9] ),
    .C(\rbzero.wall_tracer.mapY[8] ),
    .D(\rbzero.wall_tracer.mapY[10] ),
    .X(_06125_));
 sky130_fd_sc_hd__inv_2 _12950_ (.A(\rbzero.wall_tracer.mapX[5] ),
    .Y(_06126_));
 sky130_fd_sc_hd__or4_1 _12951_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(\rbzero.wall_tracer.mapX[8] ),
    .C(\rbzero.wall_tracer.mapX[10] ),
    .D(\rbzero.wall_tracer.mapY[7] ),
    .X(_06127_));
 sky130_fd_sc_hd__a2111o_1 _12952_ (.A1(\rbzero.debug_overlay.playerX[5] ),
    .A2(_06126_),
    .B1(\rbzero.wall_tracer.mapX[7] ),
    .C1(\rbzero.wall_tracer.mapX[6] ),
    .D1(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__clkinv_2 _12953_ (.A(\rbzero.map_rom.i_col[4] ),
    .Y(_06129_));
 sky130_fd_sc_hd__clkinv_2 _12954_ (.A(\rbzero.map_rom.d6 ),
    .Y(_06130_));
 sky130_fd_sc_hd__o22ai_1 _12955_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_06129_),
    .B1(_06130_),
    .B2(\rbzero.debug_overlay.playerY[0] ),
    .Y(_06131_));
 sky130_fd_sc_hd__a221o_1 _12956_ (.A1(\rbzero.debug_overlay.playerY[2] ),
    .A2(_06086_),
    .B1(\rbzero.map_rom.a6 ),
    .B2(_04667_),
    .C1(_06131_),
    .X(_06132_));
 sky130_fd_sc_hd__inv_2 _12957_ (.A(\rbzero.debug_overlay.playerX[5] ),
    .Y(_06133_));
 sky130_fd_sc_hd__a22o_1 _12958_ (.A1(_04674_),
    .A2(\rbzero.map_rom.f2 ),
    .B1(\rbzero.wall_tracer.mapX[5] ),
    .B2(_06133_),
    .X(_06134_));
 sky130_fd_sc_hd__a221o_1 _12959_ (.A1(\rbzero.debug_overlay.playerX[4] ),
    .A2(_06129_),
    .B1(_06130_),
    .B2(\rbzero.debug_overlay.playerY[0] ),
    .C1(_06134_),
    .X(_06135_));
 sky130_fd_sc_hd__or4_1 _12960_ (.A(_06125_),
    .B(_06128_),
    .C(_06132_),
    .D(_06135_),
    .X(_06136_));
 sky130_fd_sc_hd__nor2_1 _12961_ (.A(_06124_),
    .B(_06136_),
    .Y(_06137_));
 sky130_fd_sc_hd__or4_1 _12962_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(\rbzero.wall_tracer.visualWallDist[6] ),
    .C(\rbzero.wall_tracer.visualWallDist[5] ),
    .D(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_06138_));
 sky130_fd_sc_hd__or4_1 _12963_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(\rbzero.wall_tracer.visualWallDist[2] ),
    .C(\rbzero.wall_tracer.visualWallDist[1] ),
    .D(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_06139_));
 sky130_fd_sc_hd__or4_1 _12964_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(\rbzero.wall_tracer.visualWallDist[-2] ),
    .C(\rbzero.wall_tracer.visualWallDist[-3] ),
    .D(_06139_),
    .X(_06140_));
 sky130_fd_sc_hd__or4_1 _12965_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(\rbzero.wall_tracer.visualWallDist[8] ),
    .C(_06138_),
    .D(_06140_),
    .X(_06141_));
 sky130_fd_sc_hd__or3b_4 _12966_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_06137_),
    .C_N(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__a22o_1 _12967_ (.A1(\rbzero.map_overlay.i_mapdx[2] ),
    .A2(_06120_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .B2(_04720_),
    .X(_06143_));
 sky130_fd_sc_hd__clkbuf_4 _12968_ (.A(\rbzero.map_rom.f4 ),
    .X(_06144_));
 sky130_fd_sc_hd__and2_1 _12969_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_06144_),
    .X(_06145_));
 sky130_fd_sc_hd__nor2_1 _12970_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_06144_),
    .Y(_06146_));
 sky130_fd_sc_hd__xnor2_1 _12971_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(\rbzero.map_rom.f1 ),
    .Y(_06147_));
 sky130_fd_sc_hd__o221a_1 _12972_ (.A1(\rbzero.map_overlay.i_mapdx[1] ),
    .A2(_06117_),
    .B1(_06120_),
    .B2(\rbzero.map_overlay.i_mapdx[2] ),
    .C1(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__o221a_1 _12973_ (.A1(_04721_),
    .A2(_06113_),
    .B1(_06145_),
    .B2(_06146_),
    .C1(_06148_),
    .X(_06149_));
 sky130_fd_sc_hd__a21o_1 _12974_ (.A1(_04720_),
    .A2(_04725_),
    .B1(\rbzero.map_rom.i_col[4] ),
    .X(_06150_));
 sky130_fd_sc_hd__and4bb_2 _12975_ (.A_N(_06142_),
    .B_N(_06143_),
    .C(_06149_),
    .D(_06150_),
    .X(_06151_));
 sky130_fd_sc_hd__xor2_1 _12976_ (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .B(\rbzero.map_rom.b6 ),
    .X(_06152_));
 sky130_fd_sc_hd__a221o_1 _12977_ (.A1(\rbzero.map_overlay.i_mapdy[1] ),
    .A2(_06089_),
    .B1(_06121_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__xnor2_1 _12978_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(\rbzero.map_rom.a6 ),
    .Y(_06154_));
 sky130_fd_sc_hd__o221a_1 _12979_ (.A1(_04738_),
    .A2(_06088_),
    .B1(_06121_),
    .B2(\rbzero.map_overlay.i_mapdy[4] ),
    .C1(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__o221a_1 _12980_ (.A1(\rbzero.map_overlay.i_mapdy[0] ),
    .A2(_06130_),
    .B1(_06089_),
    .B2(\rbzero.map_overlay.i_mapdy[1] ),
    .C1(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__or2_1 _12981_ (.A(_06088_),
    .B(\rbzero.map_rom.c6 ),
    .X(_06157_));
 sky130_fd_sc_hd__or4_1 _12982_ (.A(\rbzero.map_rom.b6 ),
    .B(\rbzero.map_rom.a6 ),
    .C(\rbzero.map_rom.i_row[4] ),
    .D(_06157_),
    .X(_06158_));
 sky130_fd_sc_hd__and4bb_2 _12983_ (.A_N(_06142_),
    .B_N(_06153_),
    .C(_06156_),
    .D(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__nor2_2 _12984_ (.A(_06151_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__nand2_2 _12985_ (.A(_06106_),
    .B(_06160_),
    .Y(_06161_));
 sky130_fd_sc_hd__inv_2 _12986_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .Y(_06162_));
 sky130_fd_sc_hd__or2_1 _12987_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(_06162_),
    .X(_06163_));
 sky130_fd_sc_hd__inv_2 _12988_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .Y(_06164_));
 sky130_fd_sc_hd__inv_2 _12989_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .Y(_06165_));
 sky130_fd_sc_hd__a22o_1 _12990_ (.A1(\rbzero.wall_tracer.trackDistY[9] ),
    .A2(_06162_),
    .B1(\rbzero.wall_tracer.trackDistY[8] ),
    .B2(_06165_),
    .X(_06166_));
 sky130_fd_sc_hd__inv_2 _12991_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .Y(_06167_));
 sky130_fd_sc_hd__inv_2 _12992_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .Y(_06168_));
 sky130_fd_sc_hd__inv_2 _12993_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .Y(_06169_));
 sky130_fd_sc_hd__inv_2 _12994_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .Y(_06170_));
 sky130_fd_sc_hd__inv_2 _12995_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .Y(_06171_));
 sky130_fd_sc_hd__inv_2 _12996_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .Y(_06172_));
 sky130_fd_sc_hd__inv_2 _12997_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .Y(_06173_));
 sky130_fd_sc_hd__nor2_1 _12998_ (.A(_06173_),
    .B(\rbzero.wall_tracer.trackDistX[-1] ),
    .Y(_06174_));
 sky130_fd_sc_hd__inv_2 _12999_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .Y(_06175_));
 sky130_fd_sc_hd__a22o_1 _13000_ (.A1(_06175_),
    .A2(\rbzero.wall_tracer.trackDistX[0] ),
    .B1(_06173_),
    .B2(\rbzero.wall_tracer.trackDistX[-1] ),
    .X(_06176_));
 sky130_fd_sc_hd__or2_1 _13001_ (.A(_06175_),
    .B(\rbzero.wall_tracer.trackDistX[0] ),
    .X(_06177_));
 sky130_fd_sc_hd__or3b_1 _13002_ (.A(_06174_),
    .B(_06176_),
    .C_N(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__inv_2 _13003_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .Y(_06179_));
 sky130_fd_sc_hd__inv_2 _13004_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .Y(_06180_));
 sky130_fd_sc_hd__a22o_1 _13005_ (.A1(_06179_),
    .A2(\rbzero.wall_tracer.trackDistX[-2] ),
    .B1(\rbzero.wall_tracer.trackDistX[-3] ),
    .B2(_06180_),
    .X(_06181_));
 sky130_fd_sc_hd__inv_2 _13006_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .Y(_06182_));
 sky130_fd_sc_hd__inv_2 _13007_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .Y(_06183_));
 sky130_fd_sc_hd__inv_2 _13008_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .Y(_06184_));
 sky130_fd_sc_hd__inv_2 _13009_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .Y(_06185_));
 sky130_fd_sc_hd__inv_2 _13010_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .Y(_06186_));
 sky130_fd_sc_hd__inv_2 _13011_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .Y(_06187_));
 sky130_fd_sc_hd__inv_2 _13012_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .Y(_06188_));
 sky130_fd_sc_hd__inv_2 _13013_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .Y(_06189_));
 sky130_fd_sc_hd__o211a_1 _13014_ (.A1(\rbzero.wall_tracer.trackDistY[-10] ),
    .A2(_06188_),
    .B1(\rbzero.wall_tracer.trackDistY[-11] ),
    .C1(_06189_),
    .X(_06190_));
 sky130_fd_sc_hd__a221o_1 _13015_ (.A1(\rbzero.wall_tracer.trackDistY[-9] ),
    .A2(_06187_),
    .B1(\rbzero.wall_tracer.trackDistY[-10] ),
    .B2(_06188_),
    .C1(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__o221a_1 _13016_ (.A1(\rbzero.wall_tracer.trackDistY[-8] ),
    .A2(_06186_),
    .B1(\rbzero.wall_tracer.trackDistY[-9] ),
    .B2(_06187_),
    .C1(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__a221o_1 _13017_ (.A1(_06185_),
    .A2(\rbzero.wall_tracer.trackDistY[-7] ),
    .B1(\rbzero.wall_tracer.trackDistY[-8] ),
    .B2(_06186_),
    .C1(_06192_),
    .X(_06193_));
 sky130_fd_sc_hd__o221a_1 _13018_ (.A1(\rbzero.wall_tracer.trackDistY[-6] ),
    .A2(_06184_),
    .B1(_06185_),
    .B2(\rbzero.wall_tracer.trackDistY[-7] ),
    .C1(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__a221o_1 _13019_ (.A1(\rbzero.wall_tracer.trackDistY[-5] ),
    .A2(_06183_),
    .B1(\rbzero.wall_tracer.trackDistY[-6] ),
    .B2(_06184_),
    .C1(_06194_),
    .X(_06195_));
 sky130_fd_sc_hd__o221a_1 _13020_ (.A1(\rbzero.wall_tracer.trackDistY[-4] ),
    .A2(_06182_),
    .B1(\rbzero.wall_tracer.trackDistY[-5] ),
    .B2(_06183_),
    .C1(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__inv_2 _13021_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .Y(_06197_));
 sky130_fd_sc_hd__or2_1 _13022_ (.A(_06179_),
    .B(\rbzero.wall_tracer.trackDistX[-2] ),
    .X(_06198_));
 sky130_fd_sc_hd__inv_2 _13023_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .Y(_06199_));
 sky130_fd_sc_hd__o22a_1 _13024_ (.A1(\rbzero.wall_tracer.trackDistX[1] ),
    .A2(_06199_),
    .B1(\rbzero.wall_tracer.trackDistX[-3] ),
    .B2(_06180_),
    .X(_06200_));
 sky130_fd_sc_hd__o211ai_1 _13025_ (.A1(_06197_),
    .A2(\rbzero.wall_tracer.trackDistX[-4] ),
    .B1(_06198_),
    .C1(_06200_),
    .Y(_06201_));
 sky130_fd_sc_hd__inv_2 _13026_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .Y(_06202_));
 sky130_fd_sc_hd__nand2_1 _13027_ (.A(_06181_),
    .B(_06198_),
    .Y(_06203_));
 sky130_fd_sc_hd__a2bb2o_1 _13028_ (.A1_N(_06178_),
    .A2_N(_06203_),
    .B1(_06176_),
    .B2(_06177_),
    .X(_06204_));
 sky130_fd_sc_hd__o21ai_1 _13029_ (.A1(\rbzero.wall_tracer.trackDistX[1] ),
    .A2(_06199_),
    .B1(_06204_),
    .Y(_06205_));
 sky130_fd_sc_hd__o221a_1 _13030_ (.A1(\rbzero.wall_tracer.trackDistY[2] ),
    .A2(_06172_),
    .B1(_06202_),
    .B2(\rbzero.wall_tracer.trackDistY[1] ),
    .C1(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__o41a_1 _13031_ (.A1(_06178_),
    .A2(_06181_),
    .A3(_06196_),
    .A4(_06201_),
    .B1(_06206_),
    .X(_06207_));
 sky130_fd_sc_hd__a221o_1 _13032_ (.A1(\rbzero.wall_tracer.trackDistY[3] ),
    .A2(_06171_),
    .B1(\rbzero.wall_tracer.trackDistY[2] ),
    .B2(_06172_),
    .C1(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__o221a_1 _13033_ (.A1(\rbzero.wall_tracer.trackDistY[4] ),
    .A2(_06170_),
    .B1(\rbzero.wall_tracer.trackDistY[3] ),
    .B2(_06171_),
    .C1(_06208_),
    .X(_06209_));
 sky130_fd_sc_hd__a221o_1 _13034_ (.A1(_06169_),
    .A2(\rbzero.wall_tracer.trackDistY[5] ),
    .B1(\rbzero.wall_tracer.trackDistY[4] ),
    .B2(_06170_),
    .C1(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__o221a_1 _13035_ (.A1(\rbzero.wall_tracer.trackDistY[6] ),
    .A2(_06168_),
    .B1(_06169_),
    .B2(\rbzero.wall_tracer.trackDistY[5] ),
    .C1(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__a221o_1 _13036_ (.A1(\rbzero.wall_tracer.trackDistY[7] ),
    .A2(_06167_),
    .B1(\rbzero.wall_tracer.trackDistY[6] ),
    .B2(_06168_),
    .C1(_06211_),
    .X(_06212_));
 sky130_fd_sc_hd__o221a_1 _13037_ (.A1(\rbzero.wall_tracer.trackDistY[8] ),
    .A2(_06165_),
    .B1(\rbzero.wall_tracer.trackDistY[7] ),
    .B2(_06167_),
    .C1(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__or3b_1 _13038_ (.A(_06166_),
    .B(_06213_),
    .C_N(_06163_),
    .X(_06214_));
 sky130_fd_sc_hd__o21a_1 _13039_ (.A1(_06164_),
    .A2(\rbzero.wall_tracer.trackDistY[10] ),
    .B1(_06214_),
    .X(_06215_));
 sky130_fd_sc_hd__and2_1 _13040_ (.A(_06164_),
    .B(\rbzero.wall_tracer.trackDistY[10] ),
    .X(_06216_));
 sky130_fd_sc_hd__a21o_4 _13041_ (.A1(_06163_),
    .A2(_06215_),
    .B1(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__or4_1 _13042_ (.A(_06144_),
    .B(_06113_),
    .C(\rbzero.map_rom.f2 ),
    .D(\rbzero.map_rom.i_col[4] ),
    .X(_06218_));
 sky130_fd_sc_hd__a22o_1 _13043_ (.A1(_06108_),
    .A2(_06130_),
    .B1(\rbzero.map_rom.b6 ),
    .B2(\rbzero.map_rom.f2 ),
    .X(_06219_));
 sky130_fd_sc_hd__xnor2_1 _13044_ (.A(_06113_),
    .B(\rbzero.map_rom.c6 ),
    .Y(_06220_));
 sky130_fd_sc_hd__a2111o_1 _13045_ (.A1(_06120_),
    .A2(_06086_),
    .B1(\rbzero.map_rom.a6 ),
    .C1(_06219_),
    .D1(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__a221o_1 _13046_ (.A1(_06144_),
    .A2(_06088_),
    .B1(_06218_),
    .B2(_06221_),
    .C1(\rbzero.map_rom.f1 ),
    .X(_06222_));
 sky130_fd_sc_hd__nand2_1 _13047_ (.A(_06088_),
    .B(\rbzero.map_rom.c6 ),
    .Y(_06223_));
 sky130_fd_sc_hd__nand2_1 _13048_ (.A(_06157_),
    .B(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__o2bb2a_1 _13049_ (.A1_N(_06113_),
    .A2_N(_06224_),
    .B1(_06088_),
    .B2(_06144_),
    .X(_06225_));
 sky130_fd_sc_hd__or3_1 _13050_ (.A(_06120_),
    .B(_06086_),
    .C(_06225_),
    .X(_06226_));
 sky130_fd_sc_hd__or3_1 _13051_ (.A(_06086_),
    .B(_06107_),
    .C(_06121_),
    .X(_06227_));
 sky130_fd_sc_hd__inv_2 _13052_ (.A(\rbzero.map_rom.f1 ),
    .Y(_06228_));
 sky130_fd_sc_hd__nand2_1 _13053_ (.A(_06144_),
    .B(_06113_),
    .Y(_06229_));
 sky130_fd_sc_hd__or4_1 _13054_ (.A(_06120_),
    .B(_06228_),
    .C(_06129_),
    .D(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__or4_1 _13055_ (.A(\rbzero.map_rom.f4 ),
    .B(\rbzero.map_rom.f2 ),
    .C(_06088_),
    .D(\rbzero.map_rom.b6 ),
    .X(_06231_));
 sky130_fd_sc_hd__o2111a_1 _13056_ (.A1(_06223_),
    .A2(_06227_),
    .B1(_06230_),
    .C1(_06231_),
    .D1(_06158_),
    .X(_06232_));
 sky130_fd_sc_hd__and3_1 _13057_ (.A(_06222_),
    .B(_06226_),
    .C(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__inv_2 _13058_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .Y(_06234_));
 sky130_fd_sc_hd__nor2_1 _13059_ (.A(\rbzero.map_overlay.i_othery[0] ),
    .B(_06130_),
    .Y(_06235_));
 sky130_fd_sc_hd__a221o_1 _13060_ (.A1(_06234_),
    .A2(\rbzero.map_rom.i_col[4] ),
    .B1(_06086_),
    .B2(\rbzero.map_overlay.i_othery[2] ),
    .C1(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__inv_2 _13061_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .Y(_06237_));
 sky130_fd_sc_hd__a22o_1 _13062_ (.A1(\rbzero.map_overlay.i_otherx[2] ),
    .A2(_06120_),
    .B1(\rbzero.map_rom.i_row[4] ),
    .B2(_04713_),
    .X(_06238_));
 sky130_fd_sc_hd__a221o_1 _13063_ (.A1(_06237_),
    .A2(_06144_),
    .B1(_06130_),
    .B2(\rbzero.map_overlay.i_othery[0] ),
    .C1(_06238_),
    .X(_06239_));
 sky130_fd_sc_hd__a22o_1 _13064_ (.A1(\rbzero.map_overlay.i_otherx[1] ),
    .A2(_06117_),
    .B1(_06228_),
    .B2(\rbzero.map_overlay.i_otherx[3] ),
    .X(_06240_));
 sky130_fd_sc_hd__a221o_1 _13065_ (.A1(\rbzero.map_overlay.i_otherx[4] ),
    .A2(_06129_),
    .B1(_06089_),
    .B2(\rbzero.map_overlay.i_othery[1] ),
    .C1(_06240_),
    .X(_06241_));
 sky130_fd_sc_hd__nor2_1 _13066_ (.A(\rbzero.map_overlay.i_otherx[3] ),
    .B(_06228_),
    .Y(_06242_));
 sky130_fd_sc_hd__a221o_1 _13067_ (.A1(_04708_),
    .A2(_06113_),
    .B1(_06121_),
    .B2(\rbzero.map_overlay.i_othery[4] ),
    .C1(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__o22a_1 _13068_ (.A1(\rbzero.map_overlay.i_othery[2] ),
    .A2(_06086_),
    .B1(_06107_),
    .B2(\rbzero.map_overlay.i_othery[3] ),
    .X(_06244_));
 sky130_fd_sc_hd__o21ai_1 _13069_ (.A1(\rbzero.map_overlay.i_othery[1] ),
    .A2(_06089_),
    .B1(_06244_),
    .Y(_06245_));
 sky130_fd_sc_hd__a221o_1 _13070_ (.A1(\rbzero.map_overlay.i_otherx[0] ),
    .A2(_06108_),
    .B1(_06107_),
    .B2(\rbzero.map_overlay.i_othery[3] ),
    .C1(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__or4_1 _13071_ (.A(_06239_),
    .B(_06241_),
    .C(_06243_),
    .D(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__a211o_1 _13072_ (.A1(_04705_),
    .A2(\rbzero.map_rom.f2 ),
    .B1(_06236_),
    .C1(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__xnor2_1 _13073_ (.A(_06144_),
    .B(\rbzero.map_rom.b6 ),
    .Y(_06249_));
 sky130_fd_sc_hd__xnor2_1 _13074_ (.A(_06113_),
    .B(_06088_),
    .Y(_06250_));
 sky130_fd_sc_hd__a221o_1 _13075_ (.A1(_06228_),
    .A2(_06089_),
    .B1(_06107_),
    .B2(_06120_),
    .C1(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__a221o_1 _13076_ (.A1(\rbzero.map_rom.f1 ),
    .A2(\rbzero.map_rom.c6 ),
    .B1(\rbzero.map_rom.a6 ),
    .B2(\rbzero.map_rom.f2 ),
    .C1(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__and4_1 _13077_ (.A(\rbzero.map_rom.f1 ),
    .B(\rbzero.map_rom.c6 ),
    .C(\rbzero.map_rom.a6 ),
    .D(_06121_),
    .X(_06253_));
 sky130_fd_sc_hd__or4b_1 _13078_ (.A(_06113_),
    .B(\rbzero.map_rom.i_col[4] ),
    .C(_06231_),
    .D_N(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__o21ai_2 _13079_ (.A1(_06249_),
    .A2(_06252_),
    .B1(_06254_),
    .Y(_06255_));
 sky130_fd_sc_hd__inv_2 _13080_ (.A(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__a31o_2 _13081_ (.A1(_06233_),
    .A2(_06248_),
    .A3(_06256_),
    .B1(_06142_),
    .X(_06257_));
 sky130_fd_sc_hd__and2b_1 _13082_ (.A_N(_06217_),
    .B(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__and2b_1 _13083_ (.A_N(\rbzero.trace_state[3] ),
    .B(\rbzero.trace_state[2] ),
    .X(_06259_));
 sky130_fd_sc_hd__nand2_4 _13084_ (.A(\rbzero.trace_state[1] ),
    .B(_06259_),
    .Y(_06260_));
 sky130_fd_sc_hd__or2_2 _13085_ (.A(\rbzero.trace_state[0] ),
    .B(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__buf_8 _13086_ (.A(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__buf_6 _13087_ (.A(_06262_),
    .X(_06263_));
 sky130_fd_sc_hd__a21oi_2 _13088_ (.A1(_06161_),
    .A2(_06263_),
    .B1(_04432_),
    .Y(_06264_));
 sky130_fd_sc_hd__o21ai_4 _13089_ (.A1(_06161_),
    .A2(_06258_),
    .B1(_06264_),
    .Y(_06265_));
 sky130_fd_sc_hd__nor2_2 _13090_ (.A(_06105_),
    .B(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__a32o_1 _13091_ (.A1(_06101_),
    .A2(_06102_),
    .A3(_06266_),
    .B1(_06265_),
    .B2(\rbzero.wall_tracer.mapY[6] ),
    .X(_00386_));
 sky130_fd_sc_hd__xor2_1 _13092_ (.A(\rbzero.wall_tracer.mapY[7] ),
    .B(_06077_),
    .X(_06267_));
 sky130_fd_sc_hd__a21boi_1 _13093_ (.A1(\rbzero.wall_tracer.mapY[6] ),
    .A2(_06078_),
    .B1_N(_06101_),
    .Y(_06268_));
 sky130_fd_sc_hd__xnor2_1 _13094_ (.A(_06267_),
    .B(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__a22o_1 _13095_ (.A1(\rbzero.wall_tracer.mapY[7] ),
    .A2(_06265_),
    .B1(_06266_),
    .B2(_06269_),
    .X(_00387_));
 sky130_fd_sc_hd__and2_1 _13096_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .B(_06078_),
    .X(_06270_));
 sky130_fd_sc_hd__nor2_1 _13097_ (.A(\rbzero.wall_tracer.mapY[8] ),
    .B(_06078_),
    .Y(_06271_));
 sky130_fd_sc_hd__nor2_1 _13098_ (.A(_06270_),
    .B(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__o41a_1 _13099_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(\rbzero.wall_tracer.mapY[5] ),
    .A3(\rbzero.wall_tracer.mapY[7] ),
    .A4(\rbzero.wall_tracer.mapY[6] ),
    .B1(_06077_),
    .X(_06273_));
 sky130_fd_sc_hd__a31o_1 _13100_ (.A1(_06100_),
    .A2(_06099_),
    .A3(_06267_),
    .B1(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__xor2_1 _13101_ (.A(_06272_),
    .B(_06274_),
    .X(_06275_));
 sky130_fd_sc_hd__a22o_1 _13102_ (.A1(\rbzero.wall_tracer.mapY[8] ),
    .A2(_06265_),
    .B1(_06266_),
    .B2(_06275_),
    .X(_00388_));
 sky130_fd_sc_hd__a21o_1 _13103_ (.A1(_06272_),
    .A2(_06274_),
    .B1(_06270_),
    .X(_06276_));
 sky130_fd_sc_hd__xnor2_1 _13104_ (.A(\rbzero.wall_tracer.mapY[9] ),
    .B(_06078_),
    .Y(_06277_));
 sky130_fd_sc_hd__xnor2_1 _13105_ (.A(_06276_),
    .B(_06277_),
    .Y(_06278_));
 sky130_fd_sc_hd__a22o_1 _13106_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_06265_),
    .B1(_06266_),
    .B2(_06278_),
    .X(_00389_));
 sky130_fd_sc_hd__o21a_1 _13107_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_06078_),
    .B1(_06276_),
    .X(_06279_));
 sky130_fd_sc_hd__a21oi_1 _13108_ (.A1(\rbzero.wall_tracer.mapY[9] ),
    .A2(_06078_),
    .B1(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__xnor2_1 _13109_ (.A(\rbzero.wall_tracer.mapY[10] ),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand2_1 _13110_ (.A(_06078_),
    .B(_06281_),
    .Y(_06282_));
 sky130_fd_sc_hd__or2_1 _13111_ (.A(_06078_),
    .B(_06281_),
    .X(_06283_));
 sky130_fd_sc_hd__a32o_1 _13112_ (.A1(_06266_),
    .A2(_06282_),
    .A3(_06283_),
    .B1(_06265_),
    .B2(\rbzero.wall_tracer.mapY[10] ),
    .X(_00390_));
 sky130_fd_sc_hd__and2_1 _13113_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .X(_06284_));
 sky130_fd_sc_hd__nand2_1 _13114_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_06285_));
 sky130_fd_sc_hd__or2_1 _13115_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .X(_06286_));
 sky130_fd_sc_hd__nand3_1 _13116_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .C(_06286_),
    .Y(_06287_));
 sky130_fd_sc_hd__xor2_2 _13117_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_06288_));
 sky130_fd_sc_hd__nand2_1 _13118_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_06289_));
 sky130_fd_sc_hd__or2_1 _13119_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .X(_06290_));
 sky130_fd_sc_hd__nand3_1 _13120_ (.A(_06288_),
    .B(_06289_),
    .C(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__or2_1 _13121_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_06292_));
 sky130_fd_sc_hd__and2_1 _13122_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_06293_));
 sky130_fd_sc_hd__nand2_1 _13123_ (.A(\rbzero.debug_overlay.facingX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .Y(_06294_));
 sky130_fd_sc_hd__or2b_1 _13124_ (.A(_06293_),
    .B_N(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__nand2_1 _13125_ (.A(_06292_),
    .B(_06295_),
    .Y(_06296_));
 sky130_fd_sc_hd__nor2_1 _13126_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_06297_));
 sky130_fd_sc_hd__nor2_1 _13127_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06298_));
 sky130_fd_sc_hd__nand2_2 _13128_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_06299_));
 sky130_fd_sc_hd__xnor2_4 _13129_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_06300_));
 sky130_fd_sc_hd__nand2_1 _13130_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_06301_));
 sky130_fd_sc_hd__nand2_1 _13131_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_06302_));
 sky130_fd_sc_hd__o211a_1 _13132_ (.A1(_06299_),
    .A2(_06300_),
    .B1(_06301_),
    .C1(_06302_),
    .X(_06303_));
 sky130_fd_sc_hd__nand2_1 _13133_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_06304_));
 sky130_fd_sc_hd__o31ai_4 _13134_ (.A1(_06297_),
    .A2(_06298_),
    .A3(_06303_),
    .B1(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__nor2_1 _13135_ (.A(\rbzero.debug_overlay.facingX[-5] ),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_06306_));
 sky130_fd_sc_hd__nor2_1 _13136_ (.A(_06293_),
    .B(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__and2_1 _13137_ (.A(_06292_),
    .B(_06294_),
    .X(_06308_));
 sky130_fd_sc_hd__and3b_1 _13138_ (.A_N(_06291_),
    .B(_06307_),
    .C(_06308_),
    .X(_06309_));
 sky130_fd_sc_hd__a2bb2o_1 _13139_ (.A1_N(_06291_),
    .A2_N(_06296_),
    .B1(_06305_),
    .B2(_06309_),
    .X(_06310_));
 sky130_fd_sc_hd__and2_1 _13140_ (.A(\rbzero.debug_overlay.facingX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_06311_));
 sky130_fd_sc_hd__a21bo_1 _13141_ (.A1(_06311_),
    .A2(_06290_),
    .B1_N(_06289_),
    .X(_06312_));
 sky130_fd_sc_hd__nand2_1 _13142_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_06313_));
 sky130_fd_sc_hd__or2_1 _13143_ (.A(\rbzero.debug_overlay.facingX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_06314_));
 sky130_fd_sc_hd__nand2_1 _13144_ (.A(_06313_),
    .B(_06314_),
    .Y(_06315_));
 sky130_fd_sc_hd__inv_2 _13145_ (.A(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__o2111ai_1 _13146_ (.A1(_06310_),
    .A2(_06312_),
    .B1(_06316_),
    .C1(_06285_),
    .D1(_06286_),
    .Y(_06317_));
 sky130_fd_sc_hd__nand2_1 _13147_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_06318_));
 sky130_fd_sc_hd__nor2_1 _13148_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_06319_));
 sky130_fd_sc_hd__a41o_1 _13149_ (.A1(_06285_),
    .A2(_06287_),
    .A3(_06317_),
    .A4(_06318_),
    .B1(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__or2_1 _13150_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .X(_06321_));
 sky130_fd_sc_hd__o211a_4 _13151_ (.A1(_06284_),
    .A2(_06320_),
    .B1(_04443_),
    .C1(_06321_),
    .X(_06322_));
 sky130_fd_sc_hd__inv_2 _13152_ (.A(\rbzero.wall_tracer.rcp_sel[0] ),
    .Y(_06323_));
 sky130_fd_sc_hd__buf_4 _13153_ (.A(_06323_),
    .X(_06324_));
 sky130_fd_sc_hd__a31o_1 _13154_ (.A1(_05996_),
    .A2(_05998_),
    .A3(_06029_),
    .B1(_06031_),
    .X(_06325_));
 sky130_fd_sc_hd__inv_2 _13155_ (.A(\rbzero.wall_tracer.rcp_sel[2] ),
    .Y(_06326_));
 sky130_fd_sc_hd__clkbuf_4 _13156_ (.A(_06326_),
    .X(_06327_));
 sky130_fd_sc_hd__a311o_4 _13157_ (.A1(_06033_),
    .A2(_06030_),
    .A3(_06325_),
    .B1(_05995_),
    .C1(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__o211a_1 _13158_ (.A1(\rbzero.wall_tracer.visualWallDist[5] ),
    .A2(_04428_),
    .B1(_06324_),
    .C1(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__nor2_1 _13159_ (.A(_06322_),
    .B(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__or2_1 _13160_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_04428_),
    .X(_06331_));
 sky130_fd_sc_hd__a31oi_4 _13161_ (.A1(_06324_),
    .A2(_06328_),
    .A3(_06331_),
    .B1(_06322_),
    .Y(_06332_));
 sky130_fd_sc_hd__nand2_1 _13162_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_06333_));
 sky130_fd_sc_hd__nand2_1 _13163_ (.A(_06321_),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__xnor2_2 _13164_ (.A(_06320_),
    .B(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__nand2_1 _13165_ (.A(_04444_),
    .B(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__a21o_1 _13166_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_06327_),
    .B1(_04443_),
    .X(_06337_));
 sky130_fd_sc_hd__a21o_1 _13167_ (.A1(_04428_),
    .A2(_06037_),
    .B1(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__and3_1 _13168_ (.A(_06285_),
    .B(_06287_),
    .C(_06317_),
    .X(_06339_));
 sky130_fd_sc_hd__and2b_1 _13169_ (.A_N(_06319_),
    .B(_06318_),
    .X(_06340_));
 sky130_fd_sc_hd__xnor2_2 _13170_ (.A(_06339_),
    .B(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__or2_1 _13171_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_04427_),
    .X(_06342_));
 sky130_fd_sc_hd__o311a_1 _13172_ (.A1(_06327_),
    .A2(_06039_),
    .A3(_06040_),
    .B1(_06342_),
    .C1(_06323_),
    .X(_06343_));
 sky130_fd_sc_hd__a21o_1 _13173_ (.A1(_04444_),
    .A2(_06341_),
    .B1(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__a21oi_1 _13174_ (.A1(_06336_),
    .A2(_06338_),
    .B1(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand2_1 _13175_ (.A(_06289_),
    .B(_06290_),
    .Y(_06346_));
 sky130_fd_sc_hd__a32o_1 _13176_ (.A1(_06305_),
    .A2(_06307_),
    .A3(_06308_),
    .B1(_06295_),
    .B2(_06292_),
    .X(_06347_));
 sky130_fd_sc_hd__a21oi_1 _13177_ (.A1(_06288_),
    .A2(_06347_),
    .B1(_06311_),
    .Y(_06348_));
 sky130_fd_sc_hd__xnor2_1 _13178_ (.A(_06346_),
    .B(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__nand2_1 _13179_ (.A(_04443_),
    .B(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__a21o_1 _13180_ (.A1(\rbzero.wall_tracer.visualWallDist[-2] ),
    .A2(_06327_),
    .B1(_04443_),
    .X(_06351_));
 sky130_fd_sc_hd__a31o_1 _13181_ (.A1(_04427_),
    .A2(_06071_),
    .A3(_06072_),
    .B1(_06351_),
    .X(_06352_));
 sky130_fd_sc_hd__xnor2_2 _13182_ (.A(_06288_),
    .B(_06347_),
    .Y(_06353_));
 sky130_fd_sc_hd__and3_1 _13183_ (.A(_04427_),
    .B(_06048_),
    .C(_06052_),
    .X(_06354_));
 sky130_fd_sc_hd__a21o_1 _13184_ (.A1(\rbzero.wall_tracer.visualWallDist[-3] ),
    .A2(_06327_),
    .B1(_04443_),
    .X(_06355_));
 sky130_fd_sc_hd__o2bb2a_4 _13185_ (.A1_N(_04443_),
    .A2_N(_06353_),
    .B1(_06354_),
    .B2(_06355_),
    .X(_06356_));
 sky130_fd_sc_hd__a21o_1 _13186_ (.A1(_06305_),
    .A2(_06307_),
    .B1(_06293_),
    .X(_06357_));
 sky130_fd_sc_hd__xnor2_1 _13187_ (.A(_06308_),
    .B(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__nand2_1 _13188_ (.A(_04443_),
    .B(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__a21o_1 _13189_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_06327_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06360_));
 sky130_fd_sc_hd__a21o_1 _13190_ (.A1(_04427_),
    .A2(_06056_),
    .B1(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__xnor2_1 _13191_ (.A(_06305_),
    .B(_06307_),
    .Y(_06362_));
 sky130_fd_sc_hd__a21o_1 _13192_ (.A1(\rbzero.wall_tracer.visualWallDist[-5] ),
    .A2(_06327_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06363_));
 sky130_fd_sc_hd__and3_1 _13193_ (.A(_04427_),
    .B(_06046_),
    .C(_06057_),
    .X(_06364_));
 sky130_fd_sc_hd__o2bb2a_1 _13194_ (.A1_N(\rbzero.wall_tracer.rcp_sel[0] ),
    .A2_N(_06362_),
    .B1(_06363_),
    .B2(_06364_),
    .X(_06365_));
 sky130_fd_sc_hd__xor2_4 _13195_ (.A(_06299_),
    .B(_06300_),
    .X(_06366_));
 sky130_fd_sc_hd__or2_1 _13196_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06367_));
 sky130_fd_sc_hd__o211a_1 _13197_ (.A1(_06326_),
    .A2(_06065_),
    .B1(_06367_),
    .C1(_06323_),
    .X(_06368_));
 sky130_fd_sc_hd__mux2_1 _13198_ (.A0(\rbzero.wall_tracer.visualWallDist[-11] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06369_));
 sky130_fd_sc_hd__mux2_2 _13199_ (.A0(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A1(_06369_),
    .S(_06323_),
    .X(_06370_));
 sky130_fd_sc_hd__mux2_1 _13200_ (.A0(\rbzero.wall_tracer.visualWallDist[-10] ),
    .A1(\rbzero.wall_tracer.rayAddendY[-2] ),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06371_));
 sky130_fd_sc_hd__mux2_2 _13201_ (.A0(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A1(_06371_),
    .S(_06323_),
    .X(_06372_));
 sky130_fd_sc_hd__or2_1 _13202_ (.A(_06370_),
    .B(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__or2_1 _13203_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_06374_));
 sky130_fd_sc_hd__and2_1 _13204_ (.A(_06299_),
    .B(_06374_),
    .X(_06375_));
 sky130_fd_sc_hd__mux2_1 _13205_ (.A0(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A1(_06066_),
    .S(\rbzero.wall_tracer.rcp_sel[2] ),
    .X(_06376_));
 sky130_fd_sc_hd__mux2_4 _13206_ (.A0(_06375_),
    .A1(_06376_),
    .S(_06323_),
    .X(_06377_));
 sky130_fd_sc_hd__a2111oi_4 _13207_ (.A1(\rbzero.wall_tracer.rcp_sel[0] ),
    .A2(_06366_),
    .B1(_06368_),
    .C1(_06373_),
    .D1(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__clkinv_4 _13208_ (.A(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__o21a_1 _13209_ (.A1(_06299_),
    .A2(_06300_),
    .B1(_06302_),
    .X(_06380_));
 sky130_fd_sc_hd__and2b_1 _13210_ (.A_N(_06298_),
    .B(_06301_),
    .X(_06381_));
 sky130_fd_sc_hd__xor2_4 _13211_ (.A(_06380_),
    .B(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__a21o_1 _13212_ (.A1(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A2(_06326_),
    .B1(\rbzero.wall_tracer.rcp_sel[0] ),
    .X(_06383_));
 sky130_fd_sc_hd__a21oi_1 _13213_ (.A1(_04427_),
    .A2(_06063_),
    .B1(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__a21oi_4 _13214_ (.A1(\rbzero.wall_tracer.rcp_sel[0] ),
    .A2(_06382_),
    .B1(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__or2_1 _13215_ (.A(_06379_),
    .B(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__or2_1 _13216_ (.A(_06298_),
    .B(_06303_),
    .X(_06387_));
 sky130_fd_sc_hd__and2b_1 _13217_ (.A_N(_06297_),
    .B(_06304_),
    .X(_06388_));
 sky130_fd_sc_hd__xnor2_2 _13218_ (.A(_06387_),
    .B(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__mux2_1 _13219_ (.A0(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A1(_06062_),
    .S(_04427_),
    .X(_06390_));
 sky130_fd_sc_hd__mux2_2 _13220_ (.A0(_06389_),
    .A1(_06390_),
    .S(_06323_),
    .X(_06391_));
 sky130_fd_sc_hd__a2111o_2 _13221_ (.A1(_06359_),
    .A2(_06361_),
    .B1(_06365_),
    .C1(_06386_),
    .D1(_06391_),
    .X(_06392_));
 sky130_fd_sc_hd__a211oi_4 _13222_ (.A1(_06350_),
    .A2(_06352_),
    .B1(_06356_),
    .C1(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__o21ai_1 _13223_ (.A1(_06310_),
    .A2(_06312_),
    .B1(_06316_),
    .Y(_06394_));
 sky130_fd_sc_hd__nand2_1 _13224_ (.A(_06286_),
    .B(_06285_),
    .Y(_06395_));
 sky130_fd_sc_hd__a21oi_1 _13225_ (.A1(_06313_),
    .A2(_06394_),
    .B1(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__and3_1 _13226_ (.A(_06313_),
    .B(_06394_),
    .C(_06395_),
    .X(_06397_));
 sky130_fd_sc_hd__o21ai_1 _13227_ (.A1(_06396_),
    .A2(_06397_),
    .B1(_04444_),
    .Y(_06398_));
 sky130_fd_sc_hd__a21o_1 _13228_ (.A1(\rbzero.wall_tracer.visualWallDist[0] ),
    .A2(_06327_),
    .B1(_04443_),
    .X(_06399_));
 sky130_fd_sc_hd__a31o_1 _13229_ (.A1(_04428_),
    .A2(_06044_),
    .A3(_06045_),
    .B1(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__or3_1 _13230_ (.A(_06310_),
    .B(_06312_),
    .C(_06316_),
    .X(_06401_));
 sky130_fd_sc_hd__nand2_2 _13231_ (.A(_06394_),
    .B(_06401_),
    .Y(_06402_));
 sky130_fd_sc_hd__a21oi_1 _13232_ (.A1(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2(_06327_),
    .B1(_04443_),
    .Y(_06403_));
 sky130_fd_sc_hd__o31a_1 _13233_ (.A1(_06327_),
    .A2(_06043_),
    .A3(_06054_),
    .B1(_06403_),
    .X(_06404_));
 sky130_fd_sc_hd__a21oi_2 _13234_ (.A1(_04444_),
    .A2(_06402_),
    .B1(_06404_),
    .Y(_06405_));
 sky130_fd_sc_hd__a21oi_2 _13235_ (.A1(_06398_),
    .A2(_06400_),
    .B1(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__or2_1 _13236_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_04427_),
    .X(_06407_));
 sky130_fd_sc_hd__a31oi_4 _13237_ (.A1(_06324_),
    .A2(_06328_),
    .A3(_06407_),
    .B1(_06322_),
    .Y(_06408_));
 sky130_fd_sc_hd__and3_1 _13238_ (.A(_06393_),
    .B(_06406_),
    .C(_06408_),
    .X(_06409_));
 sky130_fd_sc_hd__or2_1 _13239_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_04428_),
    .X(_06410_));
 sky130_fd_sc_hd__a31oi_4 _13240_ (.A1(_06324_),
    .A2(_06328_),
    .A3(_06410_),
    .B1(_06322_),
    .Y(_06411_));
 sky130_fd_sc_hd__a31o_1 _13241_ (.A1(_06332_),
    .A2(_06345_),
    .A3(_06409_),
    .B1(_06411_),
    .X(_06412_));
 sky130_fd_sc_hd__xor2_2 _13242_ (.A(_06330_),
    .B(_06412_),
    .X(_06413_));
 sky130_fd_sc_hd__a31o_1 _13243_ (.A1(_06324_),
    .A2(_06328_),
    .A3(_06410_),
    .B1(_06322_),
    .X(_06414_));
 sky130_fd_sc_hd__clkbuf_4 _13244_ (.A(_06414_),
    .X(_06415_));
 sky130_fd_sc_hd__a31o_1 _13245_ (.A1(_06324_),
    .A2(_06328_),
    .A3(_06331_),
    .B1(_06322_),
    .X(_06416_));
 sky130_fd_sc_hd__a21o_1 _13246_ (.A1(_06336_),
    .A2(_06338_),
    .B1(_06344_),
    .X(_06417_));
 sky130_fd_sc_hd__nand3_1 _13247_ (.A(_06393_),
    .B(_06406_),
    .C(_06408_),
    .Y(_06418_));
 sky130_fd_sc_hd__o211a_1 _13248_ (.A1(\rbzero.wall_tracer.visualWallDist[8] ),
    .A2(_04428_),
    .B1(_06324_),
    .C1(_06328_),
    .X(_06419_));
 sky130_fd_sc_hd__or2_1 _13249_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_04428_),
    .X(_06420_));
 sky130_fd_sc_hd__a31o_1 _13250_ (.A1(_06324_),
    .A2(_06328_),
    .A3(_06420_),
    .B1(_06322_),
    .X(_06421_));
 sky130_fd_sc_hd__or2_1 _13251_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_04427_),
    .X(_06422_));
 sky130_fd_sc_hd__a31oi_4 _13252_ (.A1(_06324_),
    .A2(_06328_),
    .A3(_06422_),
    .B1(_06322_),
    .Y(_06423_));
 sky130_fd_sc_hd__nor4b_1 _13253_ (.A(_06329_),
    .B(_06419_),
    .C(_06421_),
    .D_N(_06423_),
    .Y(_06424_));
 sky130_fd_sc_hd__or4b_1 _13254_ (.A(_06416_),
    .B(_06417_),
    .C(_06418_),
    .D_N(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__o21a_1 _13255_ (.A1(_06284_),
    .A2(_06320_),
    .B1(_06321_),
    .X(_06426_));
 sky130_fd_sc_hd__or2_1 _13256_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_04428_),
    .X(_06427_));
 sky130_fd_sc_hd__a21oi_1 _13257_ (.A1(_06328_),
    .A2(_06427_),
    .B1(_04444_),
    .Y(_06428_));
 sky130_fd_sc_hd__o21ba_1 _13258_ (.A1(_06324_),
    .A2(_06426_),
    .B1_N(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__a21o_1 _13259_ (.A1(_06415_),
    .A2(_06425_),
    .B1(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__and3_1 _13260_ (.A(_06332_),
    .B(_06345_),
    .C(_06409_),
    .X(_06431_));
 sky130_fd_sc_hd__a211o_1 _13261_ (.A1(_06431_),
    .A2(_06424_),
    .B1(_06428_),
    .C1(_06411_),
    .X(_06432_));
 sky130_fd_sc_hd__inv_2 _13262_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .Y(_06433_));
 sky130_fd_sc_hd__or4_1 _13263_ (.A(_06433_),
    .B(\rbzero.wall_tracer.visualWallDist[9] ),
    .C(_04428_),
    .D(_04444_),
    .X(_06434_));
 sky130_fd_sc_hd__nor2_1 _13264_ (.A(_06425_),
    .B(_06434_),
    .Y(_06435_));
 sky130_fd_sc_hd__a21oi_4 _13265_ (.A1(_06430_),
    .A2(_06432_),
    .B1(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__or2b_1 _13266_ (.A(_06329_),
    .B_N(_06423_),
    .X(_06437_));
 sky130_fd_sc_hd__or4_1 _13267_ (.A(_06416_),
    .B(_06417_),
    .C(_06418_),
    .D(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__and3_1 _13268_ (.A(_06415_),
    .B(_06421_),
    .C(_06438_),
    .X(_06439_));
 sky130_fd_sc_hd__a21oi_1 _13269_ (.A1(_06415_),
    .A2(_06438_),
    .B1(_06421_),
    .Y(_06440_));
 sky130_fd_sc_hd__nor2_1 _13270_ (.A(_06322_),
    .B(_06419_),
    .Y(_06441_));
 sky130_fd_sc_hd__o211ai_1 _13271_ (.A1(_06421_),
    .A2(_06438_),
    .B1(_06441_),
    .C1(_06415_),
    .Y(_06442_));
 sky130_fd_sc_hd__and2_1 _13272_ (.A(_06414_),
    .B(_06421_),
    .X(_06443_));
 sky130_fd_sc_hd__a211o_1 _13273_ (.A1(_06415_),
    .A2(_06438_),
    .B1(_06441_),
    .C1(_06443_),
    .X(_06444_));
 sky130_fd_sc_hd__o211a_1 _13274_ (.A1(_06439_),
    .A2(_06440_),
    .B1(_06442_),
    .C1(_06444_),
    .X(_06445_));
 sky130_fd_sc_hd__a21oi_2 _13275_ (.A1(_06330_),
    .A2(_06431_),
    .B1(_06411_),
    .Y(_06446_));
 sky130_fd_sc_hd__xor2_1 _13276_ (.A(_06423_),
    .B(_06446_),
    .X(_06447_));
 sky130_fd_sc_hd__and4b_2 _13277_ (.A_N(_06413_),
    .B(_06436_),
    .C(_06445_),
    .D(_06447_),
    .X(_06448_));
 sky130_fd_sc_hd__a21oi_1 _13278_ (.A1(_04444_),
    .A2(_06341_),
    .B1(_06343_),
    .Y(_06449_));
 sky130_fd_sc_hd__a21oi_2 _13279_ (.A1(_06393_),
    .A2(_06406_),
    .B1(_06411_),
    .Y(_06450_));
 sky130_fd_sc_hd__xnor2_1 _13280_ (.A(_06449_),
    .B(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__and2_1 _13281_ (.A(_06398_),
    .B(_06400_),
    .X(_06452_));
 sky130_fd_sc_hd__a21o_2 _13282_ (.A1(_04444_),
    .A2(_06402_),
    .B1(_06404_),
    .X(_06453_));
 sky130_fd_sc_hd__a21o_1 _13283_ (.A1(_06453_),
    .A2(_06393_),
    .B1(_06411_),
    .X(_06454_));
 sky130_fd_sc_hd__xnor2_1 _13284_ (.A(_06452_),
    .B(_06454_),
    .Y(_06455_));
 sky130_fd_sc_hd__nand2_1 _13285_ (.A(_06336_),
    .B(_06338_),
    .Y(_06456_));
 sky130_fd_sc_hd__a31o_1 _13286_ (.A1(_06449_),
    .A2(_06393_),
    .A3(_06406_),
    .B1(_06411_),
    .X(_06457_));
 sky130_fd_sc_hd__xor2_2 _13287_ (.A(_06456_),
    .B(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__or3_2 _13288_ (.A(_06451_),
    .B(_06455_),
    .C(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__or2_2 _13289_ (.A(_06411_),
    .B(_06393_),
    .X(_06460_));
 sky130_fd_sc_hd__xnor2_2 _13290_ (.A(_06405_),
    .B(_06460_),
    .Y(_06461_));
 sky130_fd_sc_hd__a21oi_2 _13291_ (.A1(_06345_),
    .A2(_06409_),
    .B1(_06411_),
    .Y(_06462_));
 sky130_fd_sc_hd__xnor2_4 _13292_ (.A(_06332_),
    .B(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__a21o_1 _13293_ (.A1(_06414_),
    .A2(_06417_),
    .B1(_06450_),
    .X(_06464_));
 sky130_fd_sc_hd__xnor2_2 _13294_ (.A(_06408_),
    .B(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__or2_1 _13295_ (.A(_06463_),
    .B(_06465_),
    .X(_06466_));
 sky130_fd_sc_hd__nor3_4 _13296_ (.A(_06459_),
    .B(_06461_),
    .C(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__and2_1 _13297_ (.A(_06448_),
    .B(_06467_),
    .X(_06468_));
 sky130_fd_sc_hd__buf_4 _13298_ (.A(_06468_),
    .X(_06469_));
 sky130_fd_sc_hd__clkbuf_4 _13299_ (.A(_06469_),
    .X(_06470_));
 sky130_fd_sc_hd__clkinv_2 _13300_ (.A(_06365_),
    .Y(_06471_));
 sky130_fd_sc_hd__nor2_1 _13301_ (.A(_06386_),
    .B(_06391_),
    .Y(_06472_));
 sky130_fd_sc_hd__nor2_2 _13302_ (.A(_06411_),
    .B(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__xnor2_4 _13303_ (.A(_06471_),
    .B(_06473_),
    .Y(_06474_));
 sky130_fd_sc_hd__and2_2 _13304_ (.A(_06359_),
    .B(_06361_),
    .X(_06475_));
 sky130_fd_sc_hd__a21oi_4 _13305_ (.A1(_06471_),
    .A2(_06472_),
    .B1(_06411_),
    .Y(_06476_));
 sky130_fd_sc_hd__xnor2_2 _13306_ (.A(_06475_),
    .B(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__nand2_2 _13307_ (.A(_06350_),
    .B(_06352_),
    .Y(_06478_));
 sky130_fd_sc_hd__o21a_2 _13308_ (.A1(_06356_),
    .A2(_06392_),
    .B1(_06415_),
    .X(_06479_));
 sky130_fd_sc_hd__xnor2_4 _13309_ (.A(_06478_),
    .B(_06479_),
    .Y(_06480_));
 sky130_fd_sc_hd__nand2_2 _13310_ (.A(_06415_),
    .B(_06392_),
    .Y(_06481_));
 sky130_fd_sc_hd__xnor2_4 _13311_ (.A(_06356_),
    .B(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__nor2_1 _13312_ (.A(_06480_),
    .B(_06482_),
    .Y(_06483_));
 sky130_fd_sc_hd__and4_1 _13313_ (.A(_06448_),
    .B(_06467_),
    .C(_06477_),
    .D(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__and2_1 _13314_ (.A(_06474_),
    .B(_06484_),
    .X(_06485_));
 sky130_fd_sc_hd__xnor2_4 _13315_ (.A(_06453_),
    .B(_06460_),
    .Y(_06486_));
 sky130_fd_sc_hd__and3_1 _13316_ (.A(_06447_),
    .B(_06436_),
    .C(_06445_),
    .X(_06487_));
 sky130_fd_sc_hd__or2_1 _13317_ (.A(_06413_),
    .B(_06463_),
    .X(_06488_));
 sky130_fd_sc_hd__or2_1 _13318_ (.A(_06459_),
    .B(_06465_),
    .X(_06489_));
 sky130_fd_sc_hd__nor2_1 _13319_ (.A(_06488_),
    .B(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__and4_1 _13320_ (.A(_06486_),
    .B(_06487_),
    .C(_06480_),
    .D(_06490_),
    .X(_06491_));
 sky130_fd_sc_hd__xor2_1 _13321_ (.A(_06478_),
    .B(_06479_),
    .X(_06492_));
 sky130_fd_sc_hd__and4_1 _13322_ (.A(_06448_),
    .B(_06467_),
    .C(_06492_),
    .D(_06482_),
    .X(_06493_));
 sky130_fd_sc_hd__or3_2 _13323_ (.A(_06485_),
    .B(_06491_),
    .C(_06493_),
    .X(_06494_));
 sky130_fd_sc_hd__inv_2 _13324_ (.A(_06370_),
    .Y(_06495_));
 sky130_fd_sc_hd__a21o_1 _13325_ (.A1(_04444_),
    .A2(_06366_),
    .B1(_06368_),
    .X(_06496_));
 sky130_fd_sc_hd__o21a_1 _13326_ (.A1(_06373_),
    .A2(_06377_),
    .B1(_06415_),
    .X(_06497_));
 sky130_fd_sc_hd__xor2_4 _13327_ (.A(_06496_),
    .B(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__clkinv_2 _13328_ (.A(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__nand2_1 _13329_ (.A(_06373_),
    .B(_06415_),
    .Y(_06500_));
 sky130_fd_sc_hd__xor2_4 _13330_ (.A(_06377_),
    .B(_06500_),
    .X(_06501_));
 sky130_fd_sc_hd__nand2_1 _13331_ (.A(_06499_),
    .B(_06501_),
    .Y(_06502_));
 sky130_fd_sc_hd__nand2_2 _13332_ (.A(_06370_),
    .B(_06415_),
    .Y(_06503_));
 sky130_fd_sc_hd__xnor2_1 _13333_ (.A(_06372_),
    .B(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__or3_2 _13334_ (.A(_06495_),
    .B(_06502_),
    .C(_06504_),
    .X(_06505_));
 sky130_fd_sc_hd__xnor2_2 _13335_ (.A(_06423_),
    .B(_06446_),
    .Y(_06506_));
 sky130_fd_sc_hd__or4bb_2 _13336_ (.A(_06506_),
    .B(_06413_),
    .C_N(_06436_),
    .D_N(_06445_),
    .X(_06507_));
 sky130_fd_sc_hd__xor2_4 _13337_ (.A(_06475_),
    .B(_06476_),
    .X(_06508_));
 sky130_fd_sc_hd__nand2_1 _13338_ (.A(_06414_),
    .B(_06386_),
    .Y(_06509_));
 sky130_fd_sc_hd__xnor2_4 _13339_ (.A(_06391_),
    .B(_06509_),
    .Y(_06510_));
 sky130_fd_sc_hd__nand2_1 _13340_ (.A(_06379_),
    .B(_06414_),
    .Y(_06511_));
 sky130_fd_sc_hd__xnor2_4 _13341_ (.A(_06385_),
    .B(_06511_),
    .Y(_06512_));
 sky130_fd_sc_hd__or4_1 _13342_ (.A(_06474_),
    .B(_06508_),
    .C(_06510_),
    .D(_06512_),
    .X(_06513_));
 sky130_fd_sc_hd__or2_1 _13343_ (.A(_06482_),
    .B(_06513_),
    .X(_06514_));
 sky130_fd_sc_hd__or4b_4 _13344_ (.A(_06507_),
    .B(_06480_),
    .C(_06514_),
    .D_N(_06467_),
    .X(_06515_));
 sky130_fd_sc_hd__a21oi_4 _13345_ (.A1(_06379_),
    .A2(_06505_),
    .B1(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__nor2_1 _13346_ (.A(_06506_),
    .B(_06488_),
    .Y(_06517_));
 sky130_fd_sc_hd__xor2_1 _13347_ (.A(_06408_),
    .B(_06464_),
    .X(_06518_));
 sky130_fd_sc_hd__nand2_1 _13348_ (.A(_06486_),
    .B(_06492_),
    .Y(_06519_));
 sky130_fd_sc_hd__or4_2 _13349_ (.A(_06477_),
    .B(_06482_),
    .C(_06489_),
    .D(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__xor2_4 _13350_ (.A(_06372_),
    .B(_06503_),
    .X(_06521_));
 sky130_fd_sc_hd__or2_1 _13351_ (.A(_06488_),
    .B(_06489_),
    .X(_06522_));
 sky130_fd_sc_hd__or3_1 _13352_ (.A(_06482_),
    .B(_06513_),
    .C(_06519_),
    .X(_06523_));
 sky130_fd_sc_hd__or4_1 _13353_ (.A(_06502_),
    .B(_06521_),
    .C(_06522_),
    .D(_06523_),
    .X(_06524_));
 sky130_fd_sc_hd__nand2_4 _13354_ (.A(_06436_),
    .B(_06445_),
    .Y(_06525_));
 sky130_fd_sc_hd__a41oi_2 _13355_ (.A1(_06517_),
    .A2(_06518_),
    .A3(_06520_),
    .A4(_06524_),
    .B1(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__or2_1 _13356_ (.A(_06516_),
    .B(_06526_),
    .X(_06527_));
 sky130_fd_sc_hd__xnor2_1 _13357_ (.A(_06344_),
    .B(_06450_),
    .Y(_06528_));
 sky130_fd_sc_hd__o22a_1 _13358_ (.A1(_06528_),
    .A2(_06458_),
    .B1(_06459_),
    .B2(_06486_),
    .X(_06529_));
 sky130_fd_sc_hd__or3_1 _13359_ (.A(_06507_),
    .B(_06466_),
    .C(_06529_),
    .X(_06530_));
 sky130_fd_sc_hd__and2_1 _13360_ (.A(_06528_),
    .B(_06455_),
    .X(_06531_));
 sky130_fd_sc_hd__o21ai_1 _13361_ (.A1(_06458_),
    .A2(_06531_),
    .B1(_06518_),
    .Y(_06532_));
 sky130_fd_sc_hd__and4bb_1 _13362_ (.A_N(_06506_),
    .B_N(_06488_),
    .C(_06436_),
    .D(_06445_),
    .X(_06533_));
 sky130_fd_sc_hd__a21bo_1 _13363_ (.A1(_06520_),
    .A2(_06532_),
    .B1_N(_06533_),
    .X(_06534_));
 sky130_fd_sc_hd__nand2_1 _13364_ (.A(_06530_),
    .B(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__inv_2 _13365_ (.A(_06535_),
    .Y(_06536_));
 sky130_fd_sc_hd__or3_4 _13366_ (.A(_06494_),
    .B(_06527_),
    .C(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__nor2_1 _13367_ (.A(_06516_),
    .B(_06526_),
    .Y(_06538_));
 sky130_fd_sc_hd__or3_4 _13368_ (.A(_06494_),
    .B(_06538_),
    .C(_06535_),
    .X(_06539_));
 sky130_fd_sc_hd__nor2_8 _13369_ (.A(_06379_),
    .B(_06515_),
    .Y(_06540_));
 sky130_fd_sc_hd__or3_2 _13370_ (.A(_06459_),
    .B(_06507_),
    .C(_06466_),
    .X(_06541_));
 sky130_fd_sc_hd__o32ai_4 _13371_ (.A1(_06463_),
    .A2(_06507_),
    .A3(_06520_),
    .B1(_06541_),
    .B2(_06486_),
    .Y(_06542_));
 sky130_fd_sc_hd__nor2_1 _13372_ (.A(_06498_),
    .B(_06501_),
    .Y(_06543_));
 sky130_fd_sc_hd__and4bb_2 _13373_ (.A_N(_06480_),
    .B_N(_06514_),
    .C(_06448_),
    .D(_06467_),
    .X(_06544_));
 sky130_fd_sc_hd__a22o_2 _13374_ (.A1(_06474_),
    .A2(_06484_),
    .B1(_06543_),
    .B2(_06544_),
    .X(_06545_));
 sky130_fd_sc_hd__or2_1 _13375_ (.A(_06439_),
    .B(_06440_),
    .X(_06546_));
 sky130_fd_sc_hd__and2_1 _13376_ (.A(_06442_),
    .B(_06444_),
    .X(_06547_));
 sky130_fd_sc_hd__nand2_1 _13377_ (.A(_06546_),
    .B(_06547_),
    .Y(_06548_));
 sky130_fd_sc_hd__nor2_1 _13378_ (.A(_06463_),
    .B(_06518_),
    .Y(_06549_));
 sky130_fd_sc_hd__or3b_1 _13379_ (.A(_06458_),
    .B(_06465_),
    .C_N(_06531_),
    .X(_06550_));
 sky130_fd_sc_hd__o31ai_1 _13380_ (.A1(_06499_),
    .A2(_06489_),
    .A3(_06523_),
    .B1(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__o21a_1 _13381_ (.A1(_06463_),
    .A2(_06551_),
    .B1(_06448_),
    .X(_06552_));
 sky130_fd_sc_hd__a221o_1 _13382_ (.A1(_06436_),
    .A2(_06548_),
    .B1(_06448_),
    .B2(_06549_),
    .C1(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__nor4_4 _13383_ (.A(_06540_),
    .B(_06542_),
    .C(_06545_),
    .D(_06553_),
    .Y(_06554_));
 sky130_fd_sc_hd__nor2_1 _13384_ (.A(_06439_),
    .B(_06440_),
    .Y(_06555_));
 sky130_fd_sc_hd__a22o_1 _13385_ (.A1(_06430_),
    .A2(_06432_),
    .B1(_06555_),
    .B2(_06547_),
    .X(_06556_));
 sky130_fd_sc_hd__a221o_1 _13386_ (.A1(_06413_),
    .A2(_06487_),
    .B1(_06533_),
    .B2(_06465_),
    .C1(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__or3b_2 _13387_ (.A(_06493_),
    .B(_06557_),
    .C_N(_06530_),
    .X(_06558_));
 sky130_fd_sc_hd__inv_2 _13388_ (.A(_06502_),
    .Y(_06559_));
 sky130_fd_sc_hd__inv_2 _13389_ (.A(_06512_),
    .Y(_06560_));
 sky130_fd_sc_hd__or4_1 _13390_ (.A(_06474_),
    .B(_06508_),
    .C(_06510_),
    .D(_06560_),
    .X(_06561_));
 sky130_fd_sc_hd__clkinv_2 _13391_ (.A(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__and4_1 _13392_ (.A(_06448_),
    .B(_06467_),
    .C(_06483_),
    .D(_06562_),
    .X(_06563_));
 sky130_fd_sc_hd__a41o_1 _13393_ (.A1(_06370_),
    .A2(_06544_),
    .A3(_06559_),
    .A4(_06521_),
    .B1(_06563_),
    .X(_06564_));
 sky130_fd_sc_hd__nor3_2 _13394_ (.A(_06545_),
    .B(_06558_),
    .C(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__or4_4 _13395_ (.A(_06494_),
    .B(_06527_),
    .C(_06554_),
    .D(_06565_),
    .X(_06566_));
 sky130_fd_sc_hd__nor2_2 _13396_ (.A(_06486_),
    .B(_06541_),
    .Y(_06567_));
 sky130_fd_sc_hd__a31o_4 _13397_ (.A1(_06537_),
    .A2(_06539_),
    .A3(_06566_),
    .B1(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__nor3_1 _13398_ (.A(_06485_),
    .B(_06491_),
    .C(_06493_),
    .Y(_06569_));
 sky130_fd_sc_hd__or4_2 _13399_ (.A(_06540_),
    .B(_06542_),
    .C(_06545_),
    .D(_06553_),
    .X(_06570_));
 sky130_fd_sc_hd__or3_1 _13400_ (.A(_06545_),
    .B(_06558_),
    .C(_06564_),
    .X(_06571_));
 sky130_fd_sc_hd__a22o_1 _13401_ (.A1(_06569_),
    .A2(_06538_),
    .B1(_06570_),
    .B2(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__and2_1 _13402_ (.A(_06566_),
    .B(_06572_),
    .X(_06573_));
 sky130_fd_sc_hd__buf_2 _13403_ (.A(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__buf_2 _13404_ (.A(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__clkbuf_4 _13405_ (.A(_06570_),
    .X(_06576_));
 sky130_fd_sc_hd__buf_4 _13406_ (.A(_06576_),
    .X(_06577_));
 sky130_fd_sc_hd__buf_4 _13407_ (.A(_06565_),
    .X(_06578_));
 sky130_fd_sc_hd__buf_4 _13408_ (.A(_06578_),
    .X(_06579_));
 sky130_fd_sc_hd__xnor2_4 _13409_ (.A(_06577_),
    .B(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__nand2_4 _13410_ (.A(_06469_),
    .B(_06568_),
    .Y(_06581_));
 sky130_fd_sc_hd__inv_2 _13411_ (.A(_06501_),
    .Y(_06582_));
 sky130_fd_sc_hd__mux4_1 _13412_ (.A0(_06512_),
    .A1(_06582_),
    .A2(_06504_),
    .A3(_06498_),
    .S0(_06554_),
    .S1(_06578_),
    .X(_06583_));
 sky130_fd_sc_hd__xnor2_4 _13413_ (.A(_06554_),
    .B(_06578_),
    .Y(_06584_));
 sky130_fd_sc_hd__inv_2 _13414_ (.A(_06510_),
    .Y(_06585_));
 sky130_fd_sc_hd__nor4_1 _13415_ (.A(_06585_),
    .B(_06545_),
    .C(_06558_),
    .D(_06564_),
    .Y(_06586_));
 sky130_fd_sc_hd__o31a_1 _13416_ (.A1(_06545_),
    .A2(_06558_),
    .A3(_06564_),
    .B1(_06474_),
    .X(_06587_));
 sky130_fd_sc_hd__xor2_1 _13417_ (.A(_06356_),
    .B(_06481_),
    .X(_06588_));
 sky130_fd_sc_hd__clkbuf_4 _13418_ (.A(_06554_),
    .X(_06589_));
 sky130_fd_sc_hd__clkbuf_4 _13419_ (.A(_06571_),
    .X(_06590_));
 sky130_fd_sc_hd__o22a_1 _13420_ (.A1(_06588_),
    .A2(_06589_),
    .B1(_06590_),
    .B2(_06477_),
    .X(_06591_));
 sky130_fd_sc_hd__nand2_1 _13421_ (.A(_06584_),
    .B(_06591_),
    .Y(_06592_));
 sky130_fd_sc_hd__o31a_1 _13422_ (.A1(_06584_),
    .A2(_06586_),
    .A3(_06587_),
    .B1(_06592_),
    .X(_06593_));
 sky130_fd_sc_hd__nand2_2 _13423_ (.A(_06566_),
    .B(_06572_),
    .Y(_06594_));
 sky130_fd_sc_hd__clkbuf_4 _13424_ (.A(_06594_),
    .X(_06595_));
 sky130_fd_sc_hd__mux2_1 _13425_ (.A0(_06583_),
    .A1(_06593_),
    .S(_06595_),
    .X(_06596_));
 sky130_fd_sc_hd__and3_1 _13426_ (.A(_06569_),
    .B(_06538_),
    .C(_06570_),
    .X(_06597_));
 sky130_fd_sc_hd__buf_2 _13427_ (.A(_06597_),
    .X(_06598_));
 sky130_fd_sc_hd__nor2_2 _13428_ (.A(_06495_),
    .B(_06578_),
    .Y(_06599_));
 sky130_fd_sc_hd__nand2_4 _13429_ (.A(_06544_),
    .B(_06499_),
    .Y(_06600_));
 sky130_fd_sc_hd__a21o_1 _13430_ (.A1(_06598_),
    .A2(_06599_),
    .B1(_06600_),
    .X(_06601_));
 sky130_fd_sc_hd__nand2_4 _13431_ (.A(_06537_),
    .B(_06539_),
    .Y(_06602_));
 sky130_fd_sc_hd__clkbuf_4 _13432_ (.A(_06571_),
    .X(_06603_));
 sky130_fd_sc_hd__mux2_1 _13433_ (.A0(_06455_),
    .A1(_06461_),
    .S(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__mux2_1 _13434_ (.A0(_06480_),
    .A1(_06482_),
    .S(_06603_),
    .X(_06605_));
 sky130_fd_sc_hd__mux2_1 _13435_ (.A0(_06604_),
    .A1(_06605_),
    .S(_06576_),
    .X(_06606_));
 sky130_fd_sc_hd__mux2_1 _13436_ (.A0(_06463_),
    .A1(_06465_),
    .S(_06603_),
    .X(_06607_));
 sky130_fd_sc_hd__mux2_1 _13437_ (.A0(_06451_),
    .A1(_06458_),
    .S(_06565_),
    .X(_06608_));
 sky130_fd_sc_hd__mux2_1 _13438_ (.A0(_06607_),
    .A1(_06608_),
    .S(_06576_),
    .X(_06609_));
 sky130_fd_sc_hd__nand2_1 _13439_ (.A(_06569_),
    .B(_06538_),
    .Y(_06610_));
 sky130_fd_sc_hd__mux2_1 _13440_ (.A0(_06606_),
    .A1(_06609_),
    .S(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__nor2_1 _13441_ (.A(_06546_),
    .B(_06579_),
    .Y(_06612_));
 sky130_fd_sc_hd__clkbuf_4 _13442_ (.A(_06590_),
    .X(_06613_));
 sky130_fd_sc_hd__mux2_1 _13443_ (.A0(_06506_),
    .A1(_06413_),
    .S(_06613_),
    .X(_06614_));
 sky130_fd_sc_hd__mux2_1 _13444_ (.A0(_06612_),
    .A1(_06614_),
    .S(_06577_),
    .X(_06615_));
 sky130_fd_sc_hd__a211o_1 _13445_ (.A1(_06602_),
    .A2(_06611_),
    .B1(_06615_),
    .C1(_06469_),
    .X(_06616_));
 sky130_fd_sc_hd__o211ai_4 _13446_ (.A1(_06581_),
    .A2(_06596_),
    .B1(_06601_),
    .C1(_06616_),
    .Y(_06617_));
 sky130_fd_sc_hd__nor2_1 _13447_ (.A(_06494_),
    .B(_06527_),
    .Y(_06618_));
 sky130_fd_sc_hd__buf_2 _13448_ (.A(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__mux2_1 _13449_ (.A0(_06477_),
    .A1(_06588_),
    .S(_06578_),
    .X(_06620_));
 sky130_fd_sc_hd__mux2_1 _13450_ (.A0(_06486_),
    .A1(_06492_),
    .S(_06603_),
    .X(_06621_));
 sky130_fd_sc_hd__mux2_1 _13451_ (.A0(_06620_),
    .A1(_06621_),
    .S(_06554_),
    .X(_06622_));
 sky130_fd_sc_hd__and2_1 _13452_ (.A(_06619_),
    .B(_06622_),
    .X(_06623_));
 sky130_fd_sc_hd__mux2_1 _13453_ (.A0(_06451_),
    .A1(_06455_),
    .S(_06603_),
    .X(_06624_));
 sky130_fd_sc_hd__mux2_1 _13454_ (.A0(_06458_),
    .A1(_06465_),
    .S(_06578_),
    .X(_06625_));
 sky130_fd_sc_hd__mux2_1 _13455_ (.A0(_06624_),
    .A1(_06625_),
    .S(_06589_),
    .X(_06626_));
 sky130_fd_sc_hd__o21ai_1 _13456_ (.A1(_06619_),
    .A2(_06626_),
    .B1(_06602_),
    .Y(_06627_));
 sky130_fd_sc_hd__mux4_1 _13457_ (.A0(_06495_),
    .A1(_06499_),
    .A2(_06501_),
    .A3(_06521_),
    .S0(_06590_),
    .S1(_06554_),
    .X(_06628_));
 sky130_fd_sc_hd__mux4_1 _13458_ (.A0(_06474_),
    .A1(_06510_),
    .A2(_06512_),
    .A3(_06508_),
    .S0(_06590_),
    .S1(_06576_),
    .X(_06629_));
 sky130_fd_sc_hd__a21oi_1 _13459_ (.A1(_06566_),
    .A2(_06572_),
    .B1(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__a31oi_4 _13460_ (.A1(_06537_),
    .A2(_06539_),
    .A3(_06566_),
    .B1(_06567_),
    .Y(_06631_));
 sky130_fd_sc_hd__nand2_4 _13461_ (.A(_06448_),
    .B(_06467_),
    .Y(_06632_));
 sky130_fd_sc_hd__buf_4 _13462_ (.A(_06632_),
    .X(_06633_));
 sky130_fd_sc_hd__a2111o_1 _13463_ (.A1(_06574_),
    .A2(_06628_),
    .B1(_06630_),
    .C1(_06631_),
    .D1(_06633_),
    .X(_06634_));
 sky130_fd_sc_hd__mux2_1 _13464_ (.A0(_06413_),
    .A1(_06463_),
    .S(_06590_),
    .X(_06635_));
 sky130_fd_sc_hd__mux2_1 _13465_ (.A0(_06506_),
    .A1(_06555_),
    .S(_06578_),
    .X(_06636_));
 sky130_fd_sc_hd__mux2_1 _13466_ (.A0(_06635_),
    .A1(_06636_),
    .S(_06589_),
    .X(_06637_));
 sky130_fd_sc_hd__inv_2 _13467_ (.A(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__o211a_2 _13468_ (.A1(_06623_),
    .A2(_06627_),
    .B1(_06634_),
    .C1(_06638_),
    .X(_06639_));
 sky130_fd_sc_hd__buf_4 _13469_ (.A(_06639_),
    .X(_06640_));
 sky130_fd_sc_hd__clkbuf_4 _13470_ (.A(_06610_),
    .X(_06641_));
 sky130_fd_sc_hd__mux2_1 _13471_ (.A0(_06508_),
    .A1(_06482_),
    .S(_06565_),
    .X(_06642_));
 sky130_fd_sc_hd__mux2_1 _13472_ (.A0(_06474_),
    .A1(_06510_),
    .S(_06603_),
    .X(_06643_));
 sky130_fd_sc_hd__mux2_1 _13473_ (.A0(_06642_),
    .A1(_06643_),
    .S(_06570_),
    .X(_06644_));
 sky130_fd_sc_hd__nand2_1 _13474_ (.A(_06521_),
    .B(_06590_),
    .Y(_06645_));
 sky130_fd_sc_hd__o211a_1 _13475_ (.A1(_06582_),
    .A2(_06590_),
    .B1(_06598_),
    .C1(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__and3_1 _13476_ (.A(_06569_),
    .B(_06538_),
    .C(_06554_),
    .X(_06647_));
 sky130_fd_sc_hd__mux2_1 _13477_ (.A0(_06512_),
    .A1(_06498_),
    .S(_06603_),
    .X(_06648_));
 sky130_fd_sc_hd__a22o_1 _13478_ (.A1(_06537_),
    .A2(_06539_),
    .B1(_06647_),
    .B2(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__a211o_1 _13479_ (.A1(_06641_),
    .A2(_06644_),
    .B1(_06646_),
    .C1(_06649_),
    .X(_06650_));
 sky130_fd_sc_hd__nand2_1 _13480_ (.A(_06618_),
    .B(_06536_),
    .Y(_06651_));
 sky130_fd_sc_hd__mux2_1 _13481_ (.A0(_06461_),
    .A1(_06480_),
    .S(_06603_),
    .X(_06652_));
 sky130_fd_sc_hd__mux2_1 _13482_ (.A0(_06624_),
    .A1(_06652_),
    .S(_06576_),
    .X(_06653_));
 sky130_fd_sc_hd__or2_2 _13483_ (.A(_06651_),
    .B(_06653_),
    .X(_06654_));
 sky130_fd_sc_hd__nor2_8 _13484_ (.A(_06632_),
    .B(_06631_),
    .Y(_06655_));
 sky130_fd_sc_hd__o211a_1 _13485_ (.A1(_06370_),
    .A2(_06590_),
    .B1(_06645_),
    .C1(_06584_),
    .X(_06656_));
 sky130_fd_sc_hd__and2_2 _13486_ (.A(_06594_),
    .B(_06656_),
    .X(_06657_));
 sky130_fd_sc_hd__a32o_4 _13487_ (.A1(_06633_),
    .A2(_06650_),
    .A3(_06654_),
    .B1(_06655_),
    .B2(_06657_),
    .X(_06658_));
 sky130_fd_sc_hd__a21o_1 _13488_ (.A1(_06508_),
    .A2(_06578_),
    .B1(_06587_),
    .X(_06659_));
 sky130_fd_sc_hd__a211o_1 _13489_ (.A1(_06512_),
    .A2(_06590_),
    .B1(_06586_),
    .C1(_06554_),
    .X(_06660_));
 sky130_fd_sc_hd__o21a_1 _13490_ (.A1(_06576_),
    .A2(_06659_),
    .B1(_06660_),
    .X(_06661_));
 sky130_fd_sc_hd__or2_1 _13491_ (.A(_06619_),
    .B(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__nand2_1 _13492_ (.A(_06618_),
    .B(_06576_),
    .Y(_06663_));
 sky130_fd_sc_hd__nor2_1 _13493_ (.A(_06521_),
    .B(_06590_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand2_1 _13494_ (.A(_06618_),
    .B(_06589_),
    .Y(_06665_));
 sky130_fd_sc_hd__mux2_1 _13495_ (.A0(_06498_),
    .A1(_06582_),
    .S(_06603_),
    .X(_06666_));
 sky130_fd_sc_hd__o32a_1 _13496_ (.A1(_06663_),
    .A2(_06599_),
    .A3(_06664_),
    .B1(_06665_),
    .B2(_06666_),
    .X(_06667_));
 sky130_fd_sc_hd__and2_1 _13497_ (.A(_06537_),
    .B(_06539_),
    .X(_06668_));
 sky130_fd_sc_hd__clkbuf_4 _13498_ (.A(_06668_),
    .X(_06669_));
 sky130_fd_sc_hd__nor2_2 _13499_ (.A(_06469_),
    .B(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__a32o_1 _13500_ (.A1(_06662_),
    .A2(_06667_),
    .A3(_06670_),
    .B1(_06611_),
    .B2(_06525_),
    .X(_06671_));
 sky130_fd_sc_hd__mux2_1 _13501_ (.A0(_06605_),
    .A1(_06659_),
    .S(_06576_),
    .X(_06672_));
 sky130_fd_sc_hd__a21o_1 _13502_ (.A1(_06512_),
    .A2(_06603_),
    .B1(_06586_),
    .X(_06673_));
 sky130_fd_sc_hd__a22o_1 _13503_ (.A1(_06647_),
    .A2(_06673_),
    .B1(_06666_),
    .B2(_06598_),
    .X(_06674_));
 sky130_fd_sc_hd__a211o_1 _13504_ (.A1(_06641_),
    .A2(_06672_),
    .B1(_06674_),
    .C1(_06669_),
    .X(_06675_));
 sky130_fd_sc_hd__mux2_1 _13505_ (.A0(_06604_),
    .A1(_06608_),
    .S(_06554_),
    .X(_06676_));
 sky130_fd_sc_hd__or2_1 _13506_ (.A(_06641_),
    .B(_06676_),
    .X(_06677_));
 sky130_fd_sc_hd__and3_1 _13507_ (.A(_06469_),
    .B(_06568_),
    .C(_06594_),
    .X(_06678_));
 sky130_fd_sc_hd__mux2_1 _13508_ (.A0(_06582_),
    .A1(_06504_),
    .S(_06578_),
    .X(_06679_));
 sky130_fd_sc_hd__a22o_1 _13509_ (.A1(_06589_),
    .A2(_06599_),
    .B1(_06679_),
    .B2(_06584_),
    .X(_06680_));
 sky130_fd_sc_hd__a32o_4 _13510_ (.A1(_06633_),
    .A2(_06675_),
    .A3(_06677_),
    .B1(_06678_),
    .B2(_06680_),
    .X(_06681_));
 sky130_fd_sc_hd__a21o_4 _13511_ (.A1(_06658_),
    .A2(_06671_),
    .B1(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__a32o_1 _13512_ (.A1(_06641_),
    .A2(_06576_),
    .A3(_06599_),
    .B1(_06583_),
    .B2(_06594_),
    .X(_06683_));
 sky130_fd_sc_hd__o21ai_2 _13513_ (.A1(_06651_),
    .A2(_06609_),
    .B1(_06632_),
    .Y(_06684_));
 sky130_fd_sc_hd__o211a_1 _13514_ (.A1(_06576_),
    .A2(_06659_),
    .B1(_06660_),
    .C1(_06619_),
    .X(_06685_));
 sky130_fd_sc_hd__a211oi_2 _13515_ (.A1(_06641_),
    .A2(_06606_),
    .B1(_06685_),
    .C1(_06669_),
    .Y(_06686_));
 sky130_fd_sc_hd__o2bb2a_4 _13516_ (.A1_N(_06469_),
    .A2_N(_06683_),
    .B1(_06684_),
    .B2(_06686_),
    .X(_06687_));
 sky130_fd_sc_hd__a22oi_1 _13517_ (.A1(_06643_),
    .A2(_06647_),
    .B1(_06648_),
    .B2(_06598_),
    .Y(_06688_));
 sky130_fd_sc_hd__o211a_1 _13518_ (.A1(_06619_),
    .A2(_06622_),
    .B1(_06688_),
    .C1(_06602_),
    .X(_06689_));
 sky130_fd_sc_hd__nor2_1 _13519_ (.A(_06651_),
    .B(_06626_),
    .Y(_06690_));
 sky130_fd_sc_hd__or4_1 _13520_ (.A(_06632_),
    .B(_06631_),
    .C(_06574_),
    .D(_06628_),
    .X(_06691_));
 sky130_fd_sc_hd__o31a_4 _13521_ (.A1(_06469_),
    .A2(_06689_),
    .A3(_06690_),
    .B1(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__nor2_2 _13522_ (.A(_06687_),
    .B(_06692_),
    .Y(_06693_));
 sky130_fd_sc_hd__mux2_1 _13523_ (.A0(_06644_),
    .A1(_06653_),
    .S(_06641_),
    .X(_06694_));
 sky130_fd_sc_hd__mux2_1 _13524_ (.A0(_06625_),
    .A1(_06635_),
    .S(_06589_),
    .X(_06695_));
 sky130_fd_sc_hd__o22a_1 _13525_ (.A1(_06669_),
    .A2(_06694_),
    .B1(_06695_),
    .B2(_06651_),
    .X(_06696_));
 sky130_fd_sc_hd__mux4_1 _13526_ (.A0(_06585_),
    .A1(_06499_),
    .A2(_06501_),
    .A3(_06560_),
    .S0(_06554_),
    .S1(_06578_),
    .X(_06697_));
 sky130_fd_sc_hd__nand2_1 _13527_ (.A(_06595_),
    .B(_06697_),
    .Y(_06698_));
 sky130_fd_sc_hd__o211a_1 _13528_ (.A1(_06595_),
    .A2(_06656_),
    .B1(_06698_),
    .C1(_06655_),
    .X(_06699_));
 sky130_fd_sc_hd__a21o_2 _13529_ (.A1(_06633_),
    .A2(_06696_),
    .B1(_06699_),
    .X(_06700_));
 sky130_fd_sc_hd__nor2_1 _13530_ (.A(_06641_),
    .B(_06672_),
    .Y(_06701_));
 sky130_fd_sc_hd__o21ai_2 _13531_ (.A1(_06619_),
    .A2(_06676_),
    .B1(_06602_),
    .Y(_06702_));
 sky130_fd_sc_hd__a22oi_4 _13532_ (.A1(_06598_),
    .A2(_06607_),
    .B1(_06614_),
    .B2(_06647_),
    .Y(_06703_));
 sky130_fd_sc_hd__mux4_1 _13533_ (.A0(_06474_),
    .A1(_06512_),
    .A2(_06498_),
    .A3(_06510_),
    .S0(_06589_),
    .S1(_06579_),
    .X(_06704_));
 sky130_fd_sc_hd__mux2_1 _13534_ (.A0(_06680_),
    .A1(_06704_),
    .S(_06594_),
    .X(_06705_));
 sky130_fd_sc_hd__nand2_1 _13535_ (.A(_06655_),
    .B(_06705_),
    .Y(_06706_));
 sky130_fd_sc_hd__o211ai_4 _13536_ (.A1(_06701_),
    .A2(_06702_),
    .B1(_06703_),
    .C1(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__a31o_4 _13537_ (.A1(_06682_),
    .A2(_06693_),
    .A3(_06700_),
    .B1(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__or3b_1 _13538_ (.A(_06617_),
    .B(_06640_),
    .C_N(_06708_),
    .X(_06709_));
 sky130_fd_sc_hd__clkbuf_4 _13539_ (.A(_06709_),
    .X(_06710_));
 sky130_fd_sc_hd__o21ai_1 _13540_ (.A1(_06547_),
    .A2(_06579_),
    .B1(_06633_),
    .Y(_06711_));
 sky130_fd_sc_hd__a221o_1 _13541_ (.A1(_06641_),
    .A2(_06695_),
    .B1(_06636_),
    .B2(_06577_),
    .C1(_06711_),
    .X(_06712_));
 sky130_fd_sc_hd__a31o_1 _13542_ (.A1(_06619_),
    .A2(_06535_),
    .A3(_06653_),
    .B1(_06712_),
    .X(_06713_));
 sky130_fd_sc_hd__mux4_1 _13543_ (.A0(_06480_),
    .A1(_06474_),
    .A2(_06508_),
    .A3(_06482_),
    .S0(_06579_),
    .S1(_06589_),
    .X(_06714_));
 sky130_fd_sc_hd__nor2_1 _13544_ (.A(_06595_),
    .B(_06697_),
    .Y(_06715_));
 sky130_fd_sc_hd__a211o_1 _13545_ (.A1(_06595_),
    .A2(_06714_),
    .B1(_06715_),
    .C1(_06581_),
    .X(_06716_));
 sky130_fd_sc_hd__o211ai_4 _13546_ (.A1(_06657_),
    .A2(_06600_),
    .B1(_06713_),
    .C1(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__clkbuf_4 _13547_ (.A(_06717_),
    .X(_06718_));
 sky130_fd_sc_hd__xor2_4 _13548_ (.A(_06710_),
    .B(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__buf_2 _13549_ (.A(_06719_),
    .X(_06720_));
 sky130_fd_sc_hd__inv_2 _13550_ (.A(_06639_),
    .Y(_06721_));
 sky130_fd_sc_hd__buf_2 _13551_ (.A(_06617_),
    .X(_06722_));
 sky130_fd_sc_hd__inv_2 _13552_ (.A(_06722_),
    .Y(_06723_));
 sky130_fd_sc_hd__a21o_1 _13553_ (.A1(_06721_),
    .A2(_06708_),
    .B1(_06723_),
    .X(_06724_));
 sky130_fd_sc_hd__nand2_2 _13554_ (.A(_06710_),
    .B(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__buf_4 _13555_ (.A(_06692_),
    .X(_06726_));
 sky130_fd_sc_hd__xnor2_4 _13556_ (.A(_06640_),
    .B(_06708_),
    .Y(_06727_));
 sky130_fd_sc_hd__a2bb2o_4 _13557_ (.A1_N(_06686_),
    .A2_N(_06684_),
    .B1(_06683_),
    .B2(_06469_),
    .X(_06728_));
 sky130_fd_sc_hd__clkbuf_4 _13558_ (.A(_06671_),
    .X(_06729_));
 sky130_fd_sc_hd__a21oi_2 _13559_ (.A1(_06658_),
    .A2(_06729_),
    .B1(_06681_),
    .Y(_06730_));
 sky130_fd_sc_hd__or2_1 _13560_ (.A(_06687_),
    .B(_06692_),
    .X(_06731_));
 sky130_fd_sc_hd__a21oi_4 _13561_ (.A1(_06633_),
    .A2(_06696_),
    .B1(_06699_),
    .Y(_06732_));
 sky130_fd_sc_hd__o211a_2 _13562_ (.A1(_06701_),
    .A2(_06702_),
    .B1(_06703_),
    .C1(_06706_),
    .X(_06733_));
 sky130_fd_sc_hd__or4_1 _13563_ (.A(_06730_),
    .B(_06731_),
    .C(_06732_),
    .D(_06733_),
    .X(_06734_));
 sky130_fd_sc_hd__and3_1 _13564_ (.A(_06728_),
    .B(_06708_),
    .C(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__or3b_2 _13565_ (.A(_06726_),
    .B(_06727_),
    .C_N(_06735_),
    .X(_06736_));
 sky130_fd_sc_hd__clkinv_2 _13566_ (.A(_06692_),
    .Y(_06737_));
 sky130_fd_sc_hd__xnor2_4 _13567_ (.A(_06721_),
    .B(_06708_),
    .Y(_06738_));
 sky130_fd_sc_hd__a21o_1 _13568_ (.A1(_06737_),
    .A2(_06738_),
    .B1(_06735_),
    .X(_06739_));
 sky130_fd_sc_hd__nand4_2 _13569_ (.A(_06681_),
    .B(_06725_),
    .C(_06736_),
    .D(_06739_),
    .Y(_06740_));
 sky130_fd_sc_hd__xnor2_4 _13570_ (.A(_06730_),
    .B(_06726_),
    .Y(_06741_));
 sky130_fd_sc_hd__nand2_2 _13571_ (.A(_06682_),
    .B(_06693_),
    .Y(_06742_));
 sky130_fd_sc_hd__a21o_1 _13572_ (.A1(_06682_),
    .A2(_06737_),
    .B1(_06728_),
    .X(_06743_));
 sky130_fd_sc_hd__a21oi_1 _13573_ (.A1(_06742_),
    .A2(_06743_),
    .B1(_06732_),
    .Y(_06744_));
 sky130_fd_sc_hd__nand2_1 _13574_ (.A(_06707_),
    .B(_06741_),
    .Y(_06745_));
 sky130_fd_sc_hd__xnor2_1 _13575_ (.A(_06745_),
    .B(_06744_),
    .Y(_06746_));
 sky130_fd_sc_hd__and3_1 _13576_ (.A(_06682_),
    .B(_06693_),
    .C(_06700_),
    .X(_06747_));
 sky130_fd_sc_hd__clkbuf_4 _13577_ (.A(_06747_),
    .X(_06748_));
 sky130_fd_sc_hd__a21oi_1 _13578_ (.A1(_06682_),
    .A2(_06693_),
    .B1(_06700_),
    .Y(_06749_));
 sky130_fd_sc_hd__nor2_1 _13579_ (.A(_06748_),
    .B(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__nor2_1 _13580_ (.A(_06687_),
    .B(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__a32o_1 _13581_ (.A1(_06707_),
    .A2(_06741_),
    .A3(_06744_),
    .B1(_06746_),
    .B2(_06751_),
    .X(_06752_));
 sky130_fd_sc_hd__a22o_1 _13582_ (.A1(_06681_),
    .A2(_06725_),
    .B1(_06736_),
    .B2(_06739_),
    .X(_06753_));
 sky130_fd_sc_hd__a32oi_4 _13583_ (.A1(_06633_),
    .A2(_06675_),
    .A3(_06677_),
    .B1(_06678_),
    .B2(_06680_),
    .Y(_06754_));
 sky130_fd_sc_hd__nand2_2 _13584_ (.A(_06708_),
    .B(_06734_),
    .Y(_06755_));
 sky130_fd_sc_hd__or4_1 _13585_ (.A(_06754_),
    .B(_06726_),
    .C(_06727_),
    .D(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__buf_2 _13586_ (.A(_06658_),
    .X(_06757_));
 sky130_fd_sc_hd__clkbuf_4 _13587_ (.A(_06725_),
    .X(_06758_));
 sky130_fd_sc_hd__and2_2 _13588_ (.A(_06708_),
    .B(_06734_),
    .X(_06759_));
 sky130_fd_sc_hd__a22o_1 _13589_ (.A1(_06681_),
    .A2(_06738_),
    .B1(_06759_),
    .B2(_06737_),
    .X(_06760_));
 sky130_fd_sc_hd__nand4_1 _13590_ (.A(_06757_),
    .B(_06758_),
    .C(_06756_),
    .D(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__nand2_1 _13591_ (.A(_06756_),
    .B(_06761_),
    .Y(_06762_));
 sky130_fd_sc_hd__nand3_1 _13592_ (.A(_06740_),
    .B(_06752_),
    .C(_06753_),
    .Y(_06763_));
 sky130_fd_sc_hd__a21o_1 _13593_ (.A1(_06740_),
    .A2(_06753_),
    .B1(_06752_),
    .X(_06764_));
 sky130_fd_sc_hd__and3_1 _13594_ (.A(_06762_),
    .B(_06763_),
    .C(_06764_),
    .X(_06765_));
 sky130_fd_sc_hd__a31o_1 _13595_ (.A1(_06740_),
    .A2(_06752_),
    .A3(_06753_),
    .B1(_06765_),
    .X(_06766_));
 sky130_fd_sc_hd__nand2_2 _13596_ (.A(_06378_),
    .B(_06544_),
    .Y(_06767_));
 sky130_fd_sc_hd__o21ai_1 _13597_ (.A1(_06710_),
    .A2(_06718_),
    .B1(_06767_),
    .Y(_06768_));
 sky130_fd_sc_hd__clkbuf_4 _13598_ (.A(_06768_),
    .X(_06769_));
 sky130_fd_sc_hd__nor2_1 _13599_ (.A(_06754_),
    .B(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__a32oi_4 _13600_ (.A1(_06633_),
    .A2(_06650_),
    .A3(_06654_),
    .B1(_06655_),
    .B2(_06657_),
    .Y(_06771_));
 sky130_fd_sc_hd__clkbuf_4 _13601_ (.A(_06771_),
    .X(_06772_));
 sky130_fd_sc_hd__nor2_1 _13602_ (.A(_06772_),
    .B(_06719_),
    .Y(_06773_));
 sky130_fd_sc_hd__nand2_1 _13603_ (.A(_06770_),
    .B(_06773_),
    .Y(_06774_));
 sky130_fd_sc_hd__clkinv_2 _13604_ (.A(_06719_),
    .Y(_06775_));
 sky130_fd_sc_hd__nor2_1 _13605_ (.A(_06772_),
    .B(_06768_),
    .Y(_06776_));
 sky130_fd_sc_hd__and3_1 _13606_ (.A(_06729_),
    .B(_06775_),
    .C(_06776_),
    .X(_06777_));
 sky130_fd_sc_hd__a21o_1 _13607_ (.A1(_06681_),
    .A2(_06775_),
    .B1(_06776_),
    .X(_06778_));
 sky130_fd_sc_hd__and3_1 _13608_ (.A(_06774_),
    .B(_06777_),
    .C(_06778_),
    .X(_06779_));
 sky130_fd_sc_hd__a21oi_1 _13609_ (.A1(_06774_),
    .A2(_06778_),
    .B1(_06777_),
    .Y(_06780_));
 sky130_fd_sc_hd__nor2_1 _13610_ (.A(_06779_),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__nand2_1 _13611_ (.A(_06766_),
    .B(_06781_),
    .Y(_06782_));
 sky130_fd_sc_hd__a32oi_4 _13612_ (.A1(_06662_),
    .A2(_06667_),
    .A3(_06670_),
    .B1(_06611_),
    .B2(_06525_),
    .Y(_06783_));
 sky130_fd_sc_hd__or3_1 _13613_ (.A(_06771_),
    .B(_06783_),
    .C(_06754_),
    .X(_06784_));
 sky130_fd_sc_hd__nand2_2 _13614_ (.A(_06682_),
    .B(_06784_),
    .Y(_06785_));
 sky130_fd_sc_hd__nor2_1 _13615_ (.A(_06722_),
    .B(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__mux2_1 _13616_ (.A0(_06772_),
    .A1(_06729_),
    .S(_06717_),
    .X(_06787_));
 sky130_fd_sc_hd__xnor2_1 _13617_ (.A(_06786_),
    .B(_06787_),
    .Y(_06788_));
 sky130_fd_sc_hd__nor2_1 _13618_ (.A(_06640_),
    .B(_06785_),
    .Y(_06789_));
 sky130_fd_sc_hd__clkbuf_4 _13619_ (.A(_06783_),
    .X(_06790_));
 sky130_fd_sc_hd__or2_1 _13620_ (.A(_06790_),
    .B(_06717_),
    .X(_06791_));
 sky130_fd_sc_hd__xnor2_2 _13621_ (.A(_06658_),
    .B(_06783_),
    .Y(_06792_));
 sky130_fd_sc_hd__or2_1 _13622_ (.A(_06617_),
    .B(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__xor2_1 _13623_ (.A(_06791_),
    .B(_06793_),
    .X(_06794_));
 sky130_fd_sc_hd__or2_1 _13624_ (.A(_06791_),
    .B(_06793_),
    .X(_06795_));
 sky130_fd_sc_hd__a21boi_1 _13625_ (.A1(_06789_),
    .A2(_06794_),
    .B1_N(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__xnor2_1 _13626_ (.A(_06788_),
    .B(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__xnor2_2 _13627_ (.A(_06682_),
    .B(_06692_),
    .Y(_06798_));
 sky130_fd_sc_hd__nor2_1 _13628_ (.A(_06640_),
    .B(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__a21oi_1 _13629_ (.A1(_06742_),
    .A2(_06743_),
    .B1(_06733_),
    .Y(_06800_));
 sky130_fd_sc_hd__xor2_1 _13630_ (.A(_06799_),
    .B(_06800_),
    .X(_06801_));
 sky130_fd_sc_hd__xnor2_1 _13631_ (.A(_06748_),
    .B(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__xor2_1 _13632_ (.A(_06797_),
    .B(_06802_),
    .X(_06803_));
 sky130_fd_sc_hd__xor2_1 _13633_ (.A(_06789_),
    .B(_06794_),
    .X(_06804_));
 sky130_fd_sc_hd__nor2_1 _13634_ (.A(_06790_),
    .B(_06639_),
    .Y(_06805_));
 sky130_fd_sc_hd__or3b_1 _13635_ (.A(_06617_),
    .B(_06792_),
    .C_N(_06805_),
    .X(_06806_));
 sky130_fd_sc_hd__and2_2 _13636_ (.A(_06682_),
    .B(_06784_),
    .X(_06807_));
 sky130_fd_sc_hd__xnor2_4 _13637_ (.A(_06771_),
    .B(_06783_),
    .Y(_06808_));
 sky130_fd_sc_hd__a2bb2o_1 _13638_ (.A1_N(_06790_),
    .A2_N(_06617_),
    .B1(_06721_),
    .B2(_06808_),
    .X(_06809_));
 sky130_fd_sc_hd__nand4_1 _13639_ (.A(_06707_),
    .B(_06807_),
    .C(_06806_),
    .D(_06809_),
    .Y(_06810_));
 sky130_fd_sc_hd__nand2_1 _13640_ (.A(_06806_),
    .B(_06810_),
    .Y(_06811_));
 sky130_fd_sc_hd__xor2_1 _13641_ (.A(_06804_),
    .B(_06811_),
    .X(_06812_));
 sky130_fd_sc_hd__xor2_1 _13642_ (.A(_06751_),
    .B(_06746_),
    .X(_06813_));
 sky130_fd_sc_hd__nand2_1 _13643_ (.A(_06804_),
    .B(_06811_),
    .Y(_06814_));
 sky130_fd_sc_hd__a21bo_1 _13644_ (.A1(_06812_),
    .A2(_06813_),
    .B1_N(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__and2_1 _13645_ (.A(_06803_),
    .B(_06815_),
    .X(_06816_));
 sky130_fd_sc_hd__a21oi_1 _13646_ (.A1(_06763_),
    .A2(_06764_),
    .B1(_06762_),
    .Y(_06817_));
 sky130_fd_sc_hd__xor2_1 _13647_ (.A(_06803_),
    .B(_06815_),
    .X(_06818_));
 sky130_fd_sc_hd__nor3b_1 _13648_ (.A(_06765_),
    .B(_06817_),
    .C_N(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__or3b_1 _13649_ (.A(_06732_),
    .B(_06727_),
    .C_N(_06735_),
    .X(_06820_));
 sky130_fd_sc_hd__a22o_1 _13650_ (.A1(_06728_),
    .A2(_06738_),
    .B1(_06759_),
    .B2(_06700_),
    .X(_06821_));
 sky130_fd_sc_hd__nand4_1 _13651_ (.A(_06737_),
    .B(_06725_),
    .C(_06820_),
    .D(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__a22o_1 _13652_ (.A1(_06737_),
    .A2(_06725_),
    .B1(_06820_),
    .B2(_06821_),
    .X(_06823_));
 sky130_fd_sc_hd__a22o_1 _13653_ (.A1(_06799_),
    .A2(_06800_),
    .B1(_06801_),
    .B2(_06748_),
    .X(_06824_));
 sky130_fd_sc_hd__a21oi_1 _13654_ (.A1(_06822_),
    .A2(_06823_),
    .B1(_06824_),
    .Y(_06825_));
 sky130_fd_sc_hd__and3_1 _13655_ (.A(_06824_),
    .B(_06822_),
    .C(_06823_),
    .X(_06826_));
 sky130_fd_sc_hd__a211o_1 _13656_ (.A1(_06736_),
    .A2(_06740_),
    .B1(_06825_),
    .C1(_06826_),
    .X(_06827_));
 sky130_fd_sc_hd__nand2_1 _13657_ (.A(_06736_),
    .B(_06740_),
    .Y(_06828_));
 sky130_fd_sc_hd__o21bai_1 _13658_ (.A1(_06826_),
    .A2(_06825_),
    .B1_N(_06828_),
    .Y(_06829_));
 sky130_fd_sc_hd__nand2_1 _13659_ (.A(_06767_),
    .B(_06808_),
    .Y(_06830_));
 sky130_fd_sc_hd__or2_1 _13660_ (.A(_06717_),
    .B(_06785_),
    .X(_06831_));
 sky130_fd_sc_hd__xor2_1 _13661_ (.A(_06830_),
    .B(_06831_),
    .X(_06832_));
 sky130_fd_sc_hd__a2bb2o_1 _13662_ (.A1_N(_06772_),
    .A2_N(_06791_),
    .B1(_06786_),
    .B2(_06787_),
    .X(_06833_));
 sky130_fd_sc_hd__xor2_1 _13663_ (.A(_06832_),
    .B(_06833_),
    .X(_06834_));
 sky130_fd_sc_hd__nor2_1 _13664_ (.A(_06750_),
    .B(_06733_),
    .Y(_06835_));
 sky130_fd_sc_hd__a21o_1 _13665_ (.A1(_06742_),
    .A2(_06743_),
    .B1(_06640_),
    .X(_06836_));
 sky130_fd_sc_hd__nor2_1 _13666_ (.A(_06722_),
    .B(_06798_),
    .Y(_06837_));
 sky130_fd_sc_hd__xnor2_1 _13667_ (.A(_06836_),
    .B(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__xor2_1 _13668_ (.A(_06835_),
    .B(_06838_),
    .X(_06839_));
 sky130_fd_sc_hd__xnor2_1 _13669_ (.A(_06834_),
    .B(_06839_),
    .Y(_06840_));
 sky130_fd_sc_hd__or2_1 _13670_ (.A(_06788_),
    .B(_06796_),
    .X(_06841_));
 sky130_fd_sc_hd__o21a_1 _13671_ (.A1(_06797_),
    .A2(_06802_),
    .B1(_06841_),
    .X(_06842_));
 sky130_fd_sc_hd__xor2_1 _13672_ (.A(_06840_),
    .B(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__a21o_1 _13673_ (.A1(_06827_),
    .A2(_06829_),
    .B1(_06843_),
    .X(_06844_));
 sky130_fd_sc_hd__nand3_1 _13674_ (.A(_06827_),
    .B(_06843_),
    .C(_06829_),
    .Y(_06845_));
 sky130_fd_sc_hd__o211a_1 _13675_ (.A1(_06816_),
    .A2(_06819_),
    .B1(_06844_),
    .C1(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__a211oi_1 _13676_ (.A1(_06845_),
    .A2(_06844_),
    .B1(_06819_),
    .C1(_06816_),
    .Y(_06847_));
 sky130_fd_sc_hd__xnor2_1 _13677_ (.A(_06766_),
    .B(_06781_),
    .Y(_06848_));
 sky130_fd_sc_hd__or3_1 _13678_ (.A(_06846_),
    .B(_06847_),
    .C(_06848_),
    .X(_06849_));
 sky130_fd_sc_hd__or2b_1 _13679_ (.A(_06846_),
    .B_N(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__o21ai_1 _13680_ (.A1(_06840_),
    .A2(_06842_),
    .B1(_06845_),
    .Y(_06851_));
 sky130_fd_sc_hd__nor2_1 _13681_ (.A(_06830_),
    .B(_06831_),
    .Y(_06852_));
 sky130_fd_sc_hd__nor2_1 _13682_ (.A(_06785_),
    .B(_06852_),
    .Y(_06853_));
 sky130_fd_sc_hd__or2_2 _13683_ (.A(_06748_),
    .B(_06749_),
    .X(_06854_));
 sky130_fd_sc_hd__nand2_1 _13684_ (.A(_06854_),
    .B(_06721_),
    .Y(_06855_));
 sky130_fd_sc_hd__and2_1 _13685_ (.A(_06742_),
    .B(_06743_),
    .X(_06856_));
 sky130_fd_sc_hd__clkbuf_2 _13686_ (.A(_06856_),
    .X(_06857_));
 sky130_fd_sc_hd__nor2_1 _13687_ (.A(_06722_),
    .B(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__or2_1 _13688_ (.A(_06718_),
    .B(_06798_),
    .X(_06859_));
 sky130_fd_sc_hd__xnor2_1 _13689_ (.A(_06858_),
    .B(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__xnor2_2 _13690_ (.A(_06855_),
    .B(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__xnor2_2 _13691_ (.A(_06853_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__nand2_1 _13692_ (.A(_06832_),
    .B(_06833_),
    .Y(_06863_));
 sky130_fd_sc_hd__a21bo_1 _13693_ (.A1(_06834_),
    .A2(_06839_),
    .B1_N(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__xor2_2 _13694_ (.A(_06862_),
    .B(_06864_),
    .X(_06865_));
 sky130_fd_sc_hd__nand2_1 _13695_ (.A(_06820_),
    .B(_06822_),
    .Y(_06866_));
 sky130_fd_sc_hd__a22o_1 _13696_ (.A1(_06799_),
    .A2(_06858_),
    .B1(_06838_),
    .B2(_06835_),
    .X(_06867_));
 sky130_fd_sc_hd__nand2_1 _13697_ (.A(_06728_),
    .B(_06758_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand2_1 _13698_ (.A(_06700_),
    .B(_06738_),
    .Y(_06869_));
 sky130_fd_sc_hd__or2_1 _13699_ (.A(_06748_),
    .B(_06733_),
    .X(_06870_));
 sky130_fd_sc_hd__xnor2_1 _13700_ (.A(_06869_),
    .B(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__xnor2_1 _13701_ (.A(_06868_),
    .B(_06871_),
    .Y(_06872_));
 sky130_fd_sc_hd__xnor2_1 _13702_ (.A(_06867_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__xnor2_2 _13703_ (.A(_06866_),
    .B(_06873_),
    .Y(_06874_));
 sky130_fd_sc_hd__xnor2_2 _13704_ (.A(_06865_),
    .B(_06874_),
    .Y(_06875_));
 sky130_fd_sc_hd__xnor2_1 _13705_ (.A(_06851_),
    .B(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__nor2_1 _13706_ (.A(_06726_),
    .B(_06719_),
    .Y(_06877_));
 sky130_fd_sc_hd__nand2_1 _13707_ (.A(_06770_),
    .B(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__and3_1 _13708_ (.A(_06770_),
    .B(_06773_),
    .C(_06878_),
    .X(_06879_));
 sky130_fd_sc_hd__or2_1 _13709_ (.A(_06770_),
    .B(_06877_),
    .X(_06880_));
 sky130_fd_sc_hd__a21boi_1 _13710_ (.A1(_06878_),
    .A2(_06880_),
    .B1_N(_06774_),
    .Y(_06881_));
 sky130_fd_sc_hd__nor2_1 _13711_ (.A(_06879_),
    .B(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__and2b_1 _13712_ (.A_N(_06826_),
    .B(_06827_),
    .X(_06883_));
 sky130_fd_sc_hd__xnor2_1 _13713_ (.A(_06882_),
    .B(_06883_),
    .Y(_06884_));
 sky130_fd_sc_hd__xnor2_1 _13714_ (.A(_06779_),
    .B(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__xnor2_1 _13715_ (.A(_06876_),
    .B(_06885_),
    .Y(_06886_));
 sky130_fd_sc_hd__xnor2_1 _13716_ (.A(_06850_),
    .B(_06886_),
    .Y(_06887_));
 sky130_fd_sc_hd__xnor2_1 _13717_ (.A(_06782_),
    .B(_06887_),
    .Y(_06888_));
 sky130_fd_sc_hd__xnor2_1 _13718_ (.A(_06812_),
    .B(_06813_),
    .Y(_06889_));
 sky130_fd_sc_hd__a22o_1 _13719_ (.A1(_06707_),
    .A2(_06807_),
    .B1(_06806_),
    .B2(_06809_),
    .X(_06890_));
 sky130_fd_sc_hd__and3_1 _13720_ (.A(_06682_),
    .B(_06700_),
    .C(_06784_),
    .X(_06891_));
 sky130_fd_sc_hd__a21o_1 _13721_ (.A1(_06707_),
    .A2(_06808_),
    .B1(_06805_),
    .X(_06892_));
 sky130_fd_sc_hd__or4_1 _13722_ (.A(_06772_),
    .B(_06790_),
    .C(_06640_),
    .D(_06733_),
    .X(_06893_));
 sky130_fd_sc_hd__a21bo_1 _13723_ (.A1(_06891_),
    .A2(_06892_),
    .B1_N(_06893_),
    .X(_06894_));
 sky130_fd_sc_hd__and3_1 _13724_ (.A(_06810_),
    .B(_06890_),
    .C(_06894_),
    .X(_06895_));
 sky130_fd_sc_hd__a21oi_1 _13725_ (.A1(_06810_),
    .A2(_06890_),
    .B1(_06894_),
    .Y(_06896_));
 sky130_fd_sc_hd__mux2_1 _13726_ (.A0(_06726_),
    .A1(_06798_),
    .S(_06700_),
    .X(_06897_));
 sky130_fd_sc_hd__or3_1 _13727_ (.A(_06895_),
    .B(_06896_),
    .C(_06897_),
    .X(_06898_));
 sky130_fd_sc_hd__or2b_1 _13728_ (.A(_06895_),
    .B_N(_06898_),
    .X(_06899_));
 sky130_fd_sc_hd__and2b_1 _13729_ (.A_N(_06889_),
    .B(_06899_),
    .X(_06900_));
 sky130_fd_sc_hd__or4_2 _13730_ (.A(_06772_),
    .B(_06754_),
    .C(_06727_),
    .D(_06755_),
    .X(_06901_));
 sky130_fd_sc_hd__a22o_1 _13731_ (.A1(_06658_),
    .A2(_06738_),
    .B1(_06759_),
    .B2(_06681_),
    .X(_06902_));
 sky130_fd_sc_hd__nand4_2 _13732_ (.A(_06729_),
    .B(_06758_),
    .C(_06901_),
    .D(_06902_),
    .Y(_06903_));
 sky130_fd_sc_hd__a22o_1 _13733_ (.A1(_06658_),
    .A2(_06725_),
    .B1(_06756_),
    .B2(_06760_),
    .X(_06904_));
 sky130_fd_sc_hd__a21oi_1 _13734_ (.A1(_06761_),
    .A2(_06904_),
    .B1(_06748_),
    .Y(_06905_));
 sky130_fd_sc_hd__and3_1 _13735_ (.A(_06748_),
    .B(_06761_),
    .C(_06904_),
    .X(_06906_));
 sky130_fd_sc_hd__a211o_1 _13736_ (.A1(_06901_),
    .A2(_06903_),
    .B1(_06905_),
    .C1(_06906_),
    .X(_06907_));
 sky130_fd_sc_hd__xnor2_1 _13737_ (.A(_06889_),
    .B(_06899_),
    .Y(_06908_));
 sky130_fd_sc_hd__nand2_1 _13738_ (.A(_06901_),
    .B(_06903_),
    .Y(_06909_));
 sky130_fd_sc_hd__o21bai_1 _13739_ (.A1(_06906_),
    .A2(_06905_),
    .B1_N(_06909_),
    .Y(_06910_));
 sky130_fd_sc_hd__and3_1 _13740_ (.A(_06907_),
    .B(_06908_),
    .C(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__o21bai_1 _13741_ (.A1(_06765_),
    .A2(_06817_),
    .B1_N(_06818_),
    .Y(_06912_));
 sky130_fd_sc_hd__or3b_1 _13742_ (.A(_06765_),
    .B(_06817_),
    .C_N(_06818_),
    .X(_06913_));
 sky130_fd_sc_hd__o211a_1 _13743_ (.A1(_06900_),
    .A2(_06911_),
    .B1(_06912_),
    .C1(_06913_),
    .X(_06914_));
 sky130_fd_sc_hd__a211oi_1 _13744_ (.A1(_06913_),
    .A2(_06912_),
    .B1(_06911_),
    .C1(_06900_),
    .Y(_06915_));
 sky130_fd_sc_hd__a211oi_1 _13745_ (.A1(_06901_),
    .A2(_06903_),
    .B1(_06905_),
    .C1(_06906_),
    .Y(_06916_));
 sky130_fd_sc_hd__o22a_1 _13746_ (.A1(_06790_),
    .A2(_06769_),
    .B1(_06719_),
    .B2(_06772_),
    .X(_06917_));
 sky130_fd_sc_hd__nor2_1 _13747_ (.A(_06777_),
    .B(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__o21ai_2 _13748_ (.A1(_06906_),
    .A2(_06916_),
    .B1(_06918_),
    .Y(_06919_));
 sky130_fd_sc_hd__or3_1 _13749_ (.A(_06906_),
    .B(_06916_),
    .C(_06918_),
    .X(_06920_));
 sky130_fd_sc_hd__nand2_1 _13750_ (.A(_06919_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__nor3_1 _13751_ (.A(_06914_),
    .B(_06915_),
    .C(_06921_),
    .Y(_06922_));
 sky130_fd_sc_hd__o21ai_1 _13752_ (.A1(_06846_),
    .A2(_06847_),
    .B1(_06848_),
    .Y(_06923_));
 sky130_fd_sc_hd__o211a_1 _13753_ (.A1(_06914_),
    .A2(_06922_),
    .B1(_06923_),
    .C1(_06849_),
    .X(_06924_));
 sky130_fd_sc_hd__a211oi_1 _13754_ (.A1(_06849_),
    .A2(_06923_),
    .B1(_06922_),
    .C1(_06914_),
    .Y(_06925_));
 sky130_fd_sc_hd__or3_2 _13755_ (.A(_06919_),
    .B(_06924_),
    .C(_06925_),
    .X(_06926_));
 sky130_fd_sc_hd__and2b_1 _13756_ (.A_N(_06924_),
    .B(_06926_),
    .X(_06927_));
 sky130_fd_sc_hd__nor2_1 _13757_ (.A(_06888_),
    .B(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__nand2_1 _13758_ (.A(_06888_),
    .B(_06927_),
    .Y(_06929_));
 sky130_fd_sc_hd__nand2b_1 _13759_ (.A_N(_06928_),
    .B(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__o21ai_1 _13760_ (.A1(_06895_),
    .A2(_06896_),
    .B1(_06897_),
    .Y(_06931_));
 sky130_fd_sc_hd__nand2_1 _13761_ (.A(_06898_),
    .B(_06931_),
    .Y(_06932_));
 sky130_fd_sc_hd__nand3_1 _13762_ (.A(_06893_),
    .B(_06891_),
    .C(_06892_),
    .Y(_06933_));
 sky130_fd_sc_hd__a21o_1 _13763_ (.A1(_06893_),
    .A2(_06892_),
    .B1(_06891_),
    .X(_06934_));
 sky130_fd_sc_hd__nor2_1 _13764_ (.A(_06790_),
    .B(_06733_),
    .Y(_06935_));
 sky130_fd_sc_hd__nor2_1 _13765_ (.A(_06732_),
    .B(_06792_),
    .Y(_06936_));
 sky130_fd_sc_hd__nand2_1 _13766_ (.A(_06728_),
    .B(_06807_),
    .Y(_06937_));
 sky130_fd_sc_hd__xnor2_1 _13767_ (.A(_06935_),
    .B(_06936_),
    .Y(_06938_));
 sky130_fd_sc_hd__o2bb2ai_1 _13768_ (.A1_N(_06935_),
    .A2_N(_06936_),
    .B1(_06937_),
    .B2(_06938_),
    .Y(_06939_));
 sky130_fd_sc_hd__a21oi_1 _13769_ (.A1(_06933_),
    .A2(_06934_),
    .B1(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__nor2_1 _13770_ (.A(_06728_),
    .B(_06737_),
    .Y(_06941_));
 sky130_fd_sc_hd__clkbuf_4 _13771_ (.A(_06750_),
    .X(_06942_));
 sky130_fd_sc_hd__o32a_1 _13772_ (.A1(_06682_),
    .A2(_06693_),
    .A3(_06941_),
    .B1(_06942_),
    .B2(_06754_),
    .X(_06943_));
 sky130_fd_sc_hd__and3_1 _13773_ (.A(_06933_),
    .B(_06934_),
    .C(_06939_),
    .X(_06944_));
 sky130_fd_sc_hd__o21bai_1 _13774_ (.A1(_06940_),
    .A2(_06943_),
    .B1_N(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__or2b_1 _13775_ (.A(_06932_),
    .B_N(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__xnor2_1 _13776_ (.A(_06932_),
    .B(_06945_),
    .Y(_06947_));
 sky130_fd_sc_hd__a22o_1 _13777_ (.A1(_06729_),
    .A2(_06758_),
    .B1(_06901_),
    .B2(_06902_),
    .X(_06948_));
 sky130_fd_sc_hd__nand3b_1 _13778_ (.A_N(_06742_),
    .B(_06903_),
    .C(_06948_),
    .Y(_06949_));
 sky130_fd_sc_hd__a21bo_1 _13779_ (.A1(_06903_),
    .A2(_06948_),
    .B1_N(_06742_),
    .X(_06950_));
 sky130_fd_sc_hd__nor2_1 _13780_ (.A(_06790_),
    .B(_06755_),
    .Y(_06951_));
 sky130_fd_sc_hd__and3_1 _13781_ (.A(_06757_),
    .B(_06738_),
    .C(_06951_),
    .X(_06952_));
 sky130_fd_sc_hd__nand3_1 _13782_ (.A(_06949_),
    .B(_06950_),
    .C(_06952_),
    .Y(_06953_));
 sky130_fd_sc_hd__a21o_1 _13783_ (.A1(_06949_),
    .A2(_06950_),
    .B1(_06952_),
    .X(_06954_));
 sky130_fd_sc_hd__nand3_1 _13784_ (.A(_06947_),
    .B(_06953_),
    .C(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__a21oi_1 _13785_ (.A1(_06907_),
    .A2(_06910_),
    .B1(_06908_),
    .Y(_06956_));
 sky130_fd_sc_hd__a211oi_2 _13786_ (.A1(_06946_),
    .A2(_06955_),
    .B1(_06956_),
    .C1(_06911_),
    .Y(_06957_));
 sky130_fd_sc_hd__o211a_1 _13787_ (.A1(_06911_),
    .A2(_06956_),
    .B1(_06955_),
    .C1(_06946_),
    .X(_06958_));
 sky130_fd_sc_hd__clkbuf_4 _13788_ (.A(_06790_),
    .X(_06959_));
 sky130_fd_sc_hd__or2_1 _13789_ (.A(_06959_),
    .B(_06719_),
    .X(_06960_));
 sky130_fd_sc_hd__and2_1 _13790_ (.A(_06949_),
    .B(_06953_),
    .X(_06961_));
 sky130_fd_sc_hd__xnor2_1 _13791_ (.A(_06960_),
    .B(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__nor3_1 _13792_ (.A(_06957_),
    .B(_06958_),
    .C(_06962_),
    .Y(_06963_));
 sky130_fd_sc_hd__o21ai_1 _13793_ (.A1(_06914_),
    .A2(_06915_),
    .B1(_06921_),
    .Y(_06964_));
 sky130_fd_sc_hd__or3_1 _13794_ (.A(_06914_),
    .B(_06915_),
    .C(_06921_),
    .X(_06965_));
 sky130_fd_sc_hd__o211a_2 _13795_ (.A1(_06957_),
    .A2(_06963_),
    .B1(_06964_),
    .C1(_06965_),
    .X(_06966_));
 sky130_fd_sc_hd__or2_1 _13796_ (.A(_06960_),
    .B(_06961_),
    .X(_06967_));
 sky130_fd_sc_hd__a211oi_1 _13797_ (.A1(_06965_),
    .A2(_06964_),
    .B1(_06963_),
    .C1(_06957_),
    .Y(_06968_));
 sky130_fd_sc_hd__nor3_2 _13798_ (.A(_06967_),
    .B(_06966_),
    .C(_06968_),
    .Y(_06969_));
 sky130_fd_sc_hd__o21ai_2 _13799_ (.A1(_06924_),
    .A2(_06925_),
    .B1(_06919_),
    .Y(_06970_));
 sky130_fd_sc_hd__o211ai_4 _13800_ (.A1(_06966_),
    .A2(_06969_),
    .B1(_06926_),
    .C1(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__o21ai_1 _13801_ (.A1(_06966_),
    .A2(_06968_),
    .B1(_06967_),
    .Y(_06972_));
 sky130_fd_sc_hd__and2b_1 _13802_ (.A_N(_06969_),
    .B(_06972_),
    .X(_06973_));
 sky130_fd_sc_hd__nor2_1 _13803_ (.A(_06790_),
    .B(_06687_),
    .Y(_06974_));
 sky130_fd_sc_hd__nand2_1 _13804_ (.A(_06936_),
    .B(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__a22o_1 _13805_ (.A1(_06729_),
    .A2(_06700_),
    .B1(_06808_),
    .B2(_06728_),
    .X(_06976_));
 sky130_fd_sc_hd__a21bo_1 _13806_ (.A1(_06936_),
    .A2(_06974_),
    .B1_N(_06976_),
    .X(_06977_));
 sky130_fd_sc_hd__or3_1 _13807_ (.A(_06726_),
    .B(_06785_),
    .C(_06977_),
    .X(_06978_));
 sky130_fd_sc_hd__xnor2_1 _13808_ (.A(_06937_),
    .B(_06938_),
    .Y(_06979_));
 sky130_fd_sc_hd__a21oi_1 _13809_ (.A1(_06975_),
    .A2(_06978_),
    .B1(_06979_),
    .Y(_06980_));
 sky130_fd_sc_hd__nand2_1 _13810_ (.A(_06757_),
    .B(_06854_),
    .Y(_06981_));
 sky130_fd_sc_hd__nand2_2 _13811_ (.A(_06658_),
    .B(_06729_),
    .Y(_06982_));
 sky130_fd_sc_hd__or2_1 _13812_ (.A(_06982_),
    .B(_06726_),
    .X(_06983_));
 sky130_fd_sc_hd__nor2_1 _13813_ (.A(_06754_),
    .B(_06687_),
    .Y(_06984_));
 sky130_fd_sc_hd__a21oi_1 _13814_ (.A1(_06754_),
    .A2(_06983_),
    .B1(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__xnor2_1 _13815_ (.A(_06981_),
    .B(_06985_),
    .Y(_06986_));
 sky130_fd_sc_hd__and3_1 _13816_ (.A(_06979_),
    .B(_06975_),
    .C(_06978_),
    .X(_06987_));
 sky130_fd_sc_hd__nor2_1 _13817_ (.A(_06980_),
    .B(_06987_),
    .Y(_06988_));
 sky130_fd_sc_hd__and2_1 _13818_ (.A(_06986_),
    .B(_06988_),
    .X(_06989_));
 sky130_fd_sc_hd__nor2_1 _13819_ (.A(_06944_),
    .B(_06940_),
    .Y(_06990_));
 sky130_fd_sc_hd__xnor2_1 _13820_ (.A(_06990_),
    .B(_06943_),
    .Y(_06991_));
 sky130_fd_sc_hd__o21a_1 _13821_ (.A1(_06980_),
    .A2(_06989_),
    .B1(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__clkbuf_4 _13822_ (.A(_06755_),
    .X(_06993_));
 sky130_fd_sc_hd__o22a_1 _13823_ (.A1(_06790_),
    .A2(_06727_),
    .B1(_06993_),
    .B2(_06772_),
    .X(_06994_));
 sky130_fd_sc_hd__a32o_1 _13824_ (.A1(_06757_),
    .A2(_06854_),
    .A3(_06985_),
    .B1(_06681_),
    .B2(_06693_),
    .X(_06995_));
 sky130_fd_sc_hd__or3b_1 _13825_ (.A(_06952_),
    .B(_06994_),
    .C_N(_06995_),
    .X(_06996_));
 sky130_fd_sc_hd__or2_1 _13826_ (.A(_06952_),
    .B(_06994_),
    .X(_06997_));
 sky130_fd_sc_hd__or2b_1 _13827_ (.A(_06995_),
    .B_N(_06997_),
    .X(_06998_));
 sky130_fd_sc_hd__nand2_1 _13828_ (.A(_06996_),
    .B(_06998_),
    .Y(_06999_));
 sky130_fd_sc_hd__nor3_1 _13829_ (.A(_06991_),
    .B(_06980_),
    .C(_06989_),
    .Y(_07000_));
 sky130_fd_sc_hd__or3_1 _13830_ (.A(_06992_),
    .B(_06999_),
    .C(_07000_),
    .X(_07001_));
 sky130_fd_sc_hd__or2b_1 _13831_ (.A(_06992_),
    .B_N(_07001_),
    .X(_07002_));
 sky130_fd_sc_hd__a21o_1 _13832_ (.A1(_06953_),
    .A2(_06954_),
    .B1(_06947_),
    .X(_07003_));
 sky130_fd_sc_hd__and2_1 _13833_ (.A(_06955_),
    .B(_07003_),
    .X(_07004_));
 sky130_fd_sc_hd__nand2_1 _13834_ (.A(_07002_),
    .B(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__xnor2_1 _13835_ (.A(_07002_),
    .B(_07004_),
    .Y(_07006_));
 sky130_fd_sc_hd__or2_1 _13836_ (.A(_06996_),
    .B(_07006_),
    .X(_07007_));
 sky130_fd_sc_hd__o21a_1 _13837_ (.A1(_06957_),
    .A2(_06958_),
    .B1(_06962_),
    .X(_07008_));
 sky130_fd_sc_hd__a211oi_1 _13838_ (.A1(_07005_),
    .A2(_07007_),
    .B1(_06963_),
    .C1(_07008_),
    .Y(_07009_));
 sky130_fd_sc_hd__a211o_1 _13839_ (.A1(_06926_),
    .A2(_06970_),
    .B1(_06966_),
    .C1(_06969_),
    .X(_07010_));
 sky130_fd_sc_hd__nand4_1 _13840_ (.A(_06971_),
    .B(_06973_),
    .C(_07009_),
    .D(_07010_),
    .Y(_07011_));
 sky130_fd_sc_hd__a22o_1 _13841_ (.A1(_06973_),
    .A2(_07009_),
    .B1(_07010_),
    .B2(_06971_),
    .X(_07012_));
 sky130_fd_sc_hd__o211ai_1 _13842_ (.A1(_06963_),
    .A2(_07008_),
    .B1(_07005_),
    .C1(_07007_),
    .Y(_07013_));
 sky130_fd_sc_hd__and3b_1 _13843_ (.A_N(_07009_),
    .B(_07013_),
    .C(_06973_),
    .X(_07014_));
 sky130_fd_sc_hd__xor2_1 _13844_ (.A(_06996_),
    .B(_07006_),
    .X(_07015_));
 sky130_fd_sc_hd__o21ai_1 _13845_ (.A1(_06992_),
    .A2(_07000_),
    .B1(_06999_),
    .Y(_07016_));
 sky130_fd_sc_hd__nand2_1 _13846_ (.A(_07001_),
    .B(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__xnor2_1 _13847_ (.A(_06986_),
    .B(_06988_),
    .Y(_07018_));
 sky130_fd_sc_hd__nor2_1 _13848_ (.A(_06754_),
    .B(_06726_),
    .Y(_07019_));
 sky130_fd_sc_hd__nor2_1 _13849_ (.A(_06772_),
    .B(_06857_),
    .Y(_07020_));
 sky130_fd_sc_hd__xnor2_1 _13850_ (.A(_07019_),
    .B(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__nor2_1 _13851_ (.A(_06959_),
    .B(_06942_),
    .Y(_07022_));
 sky130_fd_sc_hd__xnor2_1 _13852_ (.A(_07021_),
    .B(_07022_),
    .Y(_07023_));
 sky130_fd_sc_hd__o21ai_1 _13853_ (.A1(_06726_),
    .A2(_06785_),
    .B1(_06977_),
    .Y(_07024_));
 sky130_fd_sc_hd__and2_1 _13854_ (.A(_06978_),
    .B(_07024_),
    .X(_07025_));
 sky130_fd_sc_hd__nand2_1 _13855_ (.A(_06982_),
    .B(_06681_),
    .Y(_07026_));
 sky130_fd_sc_hd__a21oi_1 _13856_ (.A1(_06737_),
    .A2(_06808_),
    .B1(_06974_),
    .Y(_07027_));
 sky130_fd_sc_hd__o22ai_2 _13857_ (.A1(_06982_),
    .A2(_06731_),
    .B1(_07026_),
    .B2(_07027_),
    .Y(_07028_));
 sky130_fd_sc_hd__xor2_1 _13858_ (.A(_07025_),
    .B(_07028_),
    .X(_07029_));
 sky130_fd_sc_hd__and3_1 _13859_ (.A(_06978_),
    .B(_07024_),
    .C(_07028_),
    .X(_07030_));
 sky130_fd_sc_hd__a21oi_1 _13860_ (.A1(_07023_),
    .A2(_07029_),
    .B1(_07030_),
    .Y(_07031_));
 sky130_fd_sc_hd__or2_1 _13861_ (.A(_07019_),
    .B(_07020_),
    .X(_07032_));
 sky130_fd_sc_hd__a32o_1 _13862_ (.A1(_06757_),
    .A2(_06728_),
    .A3(_07019_),
    .B1(_07032_),
    .B2(_07022_),
    .X(_07033_));
 sky130_fd_sc_hd__xnor2_1 _13863_ (.A(_06951_),
    .B(_07033_),
    .Y(_07034_));
 sky130_fd_sc_hd__xnor2_1 _13864_ (.A(_07018_),
    .B(_07031_),
    .Y(_07035_));
 sky130_fd_sc_hd__nor2_1 _13865_ (.A(_07034_),
    .B(_07035_),
    .Y(_07036_));
 sky130_fd_sc_hd__o21ba_1 _13866_ (.A1(_07018_),
    .A2(_07031_),
    .B1_N(_07036_),
    .X(_07037_));
 sky130_fd_sc_hd__nand2_1 _13867_ (.A(_06951_),
    .B(_07033_),
    .Y(_07038_));
 sky130_fd_sc_hd__xnor2_1 _13868_ (.A(_07017_),
    .B(_07037_),
    .Y(_07039_));
 sky130_fd_sc_hd__or2_1 _13869_ (.A(_07038_),
    .B(_07039_),
    .X(_07040_));
 sky130_fd_sc_hd__o21ai_1 _13870_ (.A1(_07017_),
    .A2(_07037_),
    .B1(_07040_),
    .Y(_07041_));
 sky130_fd_sc_hd__and2_1 _13871_ (.A(_07015_),
    .B(_07041_),
    .X(_07042_));
 sky130_fd_sc_hd__a22o_1 _13872_ (.A1(_07011_),
    .A2(_07012_),
    .B1(_07014_),
    .B2(_07042_),
    .X(_07043_));
 sky130_fd_sc_hd__xnor2_1 _13873_ (.A(_07023_),
    .B(_07029_),
    .Y(_07044_));
 sky130_fd_sc_hd__clkbuf_4 _13874_ (.A(_06798_),
    .X(_07045_));
 sky130_fd_sc_hd__o22a_1 _13875_ (.A1(_06959_),
    .A2(_06857_),
    .B1(_07045_),
    .B2(_06772_),
    .X(_07046_));
 sky130_fd_sc_hd__a211o_1 _13876_ (.A1(_07026_),
    .A2(_07027_),
    .B1(_07028_),
    .C1(_07046_),
    .X(_07047_));
 sky130_fd_sc_hd__o22a_1 _13877_ (.A1(_06728_),
    .A2(_06983_),
    .B1(_07044_),
    .B2(_07047_),
    .X(_07048_));
 sky130_fd_sc_hd__nand2_1 _13878_ (.A(_07034_),
    .B(_07035_),
    .Y(_07049_));
 sky130_fd_sc_hd__and2b_1 _13879_ (.A_N(_07036_),
    .B(_07049_),
    .X(_07050_));
 sky130_fd_sc_hd__a21oi_1 _13880_ (.A1(_06757_),
    .A2(_06729_),
    .B1(_07050_),
    .Y(_07051_));
 sky130_fd_sc_hd__a211oi_1 _13881_ (.A1(_07038_),
    .A2(_07039_),
    .B1(_07048_),
    .C1(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__o211a_1 _13882_ (.A1(_07015_),
    .A2(_07041_),
    .B1(_07052_),
    .C1(_07014_),
    .X(_07053_));
 sky130_fd_sc_hd__and4_1 _13883_ (.A(_07011_),
    .B(_07012_),
    .C(_07014_),
    .D(_07042_),
    .X(_07054_));
 sky130_fd_sc_hd__a21o_1 _13884_ (.A1(_07043_),
    .A2(_07053_),
    .B1(_07054_),
    .X(_07055_));
 sky130_fd_sc_hd__nand2_1 _13885_ (.A(_06971_),
    .B(_07011_),
    .Y(_07056_));
 sky130_fd_sc_hd__xnor2_1 _13886_ (.A(_06930_),
    .B(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__a2bb2o_1 _13887_ (.A1_N(_06930_),
    .A2_N(_07011_),
    .B1(_07055_),
    .B2(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__or2b_1 _13888_ (.A(_06883_),
    .B_N(_06882_),
    .X(_07059_));
 sky130_fd_sc_hd__a21bo_1 _13889_ (.A1(_06779_),
    .A2(_06884_),
    .B1_N(_07059_),
    .X(_07060_));
 sky130_fd_sc_hd__and2b_1 _13890_ (.A_N(_06851_),
    .B(_06875_),
    .X(_07061_));
 sky130_fd_sc_hd__and2b_1 _13891_ (.A_N(_06875_),
    .B(_06851_),
    .X(_07062_));
 sky130_fd_sc_hd__o21ba_1 _13892_ (.A1(_07061_),
    .A2(_06885_),
    .B1_N(_07062_),
    .X(_07063_));
 sky130_fd_sc_hd__or2b_1 _13893_ (.A(_06862_),
    .B_N(_06864_),
    .X(_07064_));
 sky130_fd_sc_hd__o21ai_1 _13894_ (.A1(_06865_),
    .A2(_06874_),
    .B1(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__nor2_1 _13895_ (.A(_06718_),
    .B(_06857_),
    .Y(_07066_));
 sky130_fd_sc_hd__buf_4 _13896_ (.A(_06767_),
    .X(_07067_));
 sky130_fd_sc_hd__a21oi_1 _13897_ (.A1(_07067_),
    .A2(_06741_),
    .B1(_07066_),
    .Y(_07068_));
 sky130_fd_sc_hd__a21oi_2 _13898_ (.A1(_06741_),
    .A2(_07066_),
    .B1(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__nor2_1 _13899_ (.A(_06942_),
    .B(_06722_),
    .Y(_07070_));
 sky130_fd_sc_hd__xor2_2 _13900_ (.A(_07069_),
    .B(_07070_),
    .X(_07071_));
 sky130_fd_sc_hd__a21oi_1 _13901_ (.A1(_06807_),
    .A2(_06861_),
    .B1(_06852_),
    .Y(_07072_));
 sky130_fd_sc_hd__xnor2_2 _13902_ (.A(_07071_),
    .B(_07072_),
    .Y(_07073_));
 sky130_fd_sc_hd__or2_1 _13903_ (.A(_06869_),
    .B(_06870_),
    .X(_07074_));
 sky130_fd_sc_hd__o21ai_2 _13904_ (.A1(_06868_),
    .A2(_06871_),
    .B1(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__nand2_1 _13905_ (.A(_06837_),
    .B(_07066_),
    .Y(_07076_));
 sky130_fd_sc_hd__or2b_1 _13906_ (.A(_06855_),
    .B_N(_06860_),
    .X(_07077_));
 sky130_fd_sc_hd__and2_1 _13907_ (.A(_06710_),
    .B(_06724_),
    .X(_07078_));
 sky130_fd_sc_hd__o2bb2a_1 _13908_ (.A1_N(_06748_),
    .A2_N(_06721_),
    .B1(_07078_),
    .B2(_06732_),
    .X(_07079_));
 sky130_fd_sc_hd__a31o_1 _13909_ (.A1(_06748_),
    .A2(_06721_),
    .A3(_06758_),
    .B1(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__a21oi_1 _13910_ (.A1(_07076_),
    .A2(_07077_),
    .B1(_07080_),
    .Y(_07081_));
 sky130_fd_sc_hd__and3_1 _13911_ (.A(_07076_),
    .B(_07077_),
    .C(_07080_),
    .X(_07082_));
 sky130_fd_sc_hd__nor2_1 _13912_ (.A(_07081_),
    .B(_07082_),
    .Y(_07083_));
 sky130_fd_sc_hd__xor2_2 _13913_ (.A(_07075_),
    .B(_07083_),
    .X(_07084_));
 sky130_fd_sc_hd__xor2_2 _13914_ (.A(_07073_),
    .B(_07084_),
    .X(_07085_));
 sky130_fd_sc_hd__xnor2_1 _13915_ (.A(_07065_),
    .B(_07085_),
    .Y(_07086_));
 sky130_fd_sc_hd__and2b_1 _13916_ (.A_N(_06872_),
    .B(_06867_),
    .X(_07087_));
 sky130_fd_sc_hd__a21oi_1 _13917_ (.A1(_06866_),
    .A2(_06873_),
    .B1(_07087_),
    .Y(_07088_));
 sky130_fd_sc_hd__nor2_1 _13918_ (.A(_06726_),
    .B(_06769_),
    .Y(_07089_));
 sky130_fd_sc_hd__nor2_1 _13919_ (.A(_06687_),
    .B(_06719_),
    .Y(_07090_));
 sky130_fd_sc_hd__nand2_1 _13920_ (.A(_07089_),
    .B(_07090_),
    .Y(_07091_));
 sky130_fd_sc_hd__or2_1 _13921_ (.A(_07089_),
    .B(_07090_),
    .X(_07092_));
 sky130_fd_sc_hd__and2_1 _13922_ (.A(_07091_),
    .B(_07092_),
    .X(_07093_));
 sky130_fd_sc_hd__and3_1 _13923_ (.A(_06770_),
    .B(_06877_),
    .C(_07093_),
    .X(_07094_));
 sky130_fd_sc_hd__a21oi_1 _13924_ (.A1(_06770_),
    .A2(_06877_),
    .B1(_07093_),
    .Y(_07095_));
 sky130_fd_sc_hd__nor2_1 _13925_ (.A(_07094_),
    .B(_07095_),
    .Y(_07096_));
 sky130_fd_sc_hd__xnor2_1 _13926_ (.A(_07088_),
    .B(_07096_),
    .Y(_07097_));
 sky130_fd_sc_hd__xnor2_1 _13927_ (.A(_06879_),
    .B(_07097_),
    .Y(_07098_));
 sky130_fd_sc_hd__xor2_1 _13928_ (.A(_07086_),
    .B(_07098_),
    .X(_07099_));
 sky130_fd_sc_hd__xnor2_1 _13929_ (.A(_07063_),
    .B(_07099_),
    .Y(_07100_));
 sky130_fd_sc_hd__xnor2_1 _13930_ (.A(_07060_),
    .B(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__nand2_1 _13931_ (.A(_06850_),
    .B(_06886_),
    .Y(_07102_));
 sky130_fd_sc_hd__o21a_1 _13932_ (.A1(_06782_),
    .A2(_06887_),
    .B1(_07102_),
    .X(_07103_));
 sky130_fd_sc_hd__xnor2_1 _13933_ (.A(_07101_),
    .B(_07103_),
    .Y(_07104_));
 sky130_fd_sc_hd__o21ba_1 _13934_ (.A1(_06971_),
    .A2(_06930_),
    .B1_N(_06928_),
    .X(_07105_));
 sky130_fd_sc_hd__xor2_1 _13935_ (.A(_07104_),
    .B(_07105_),
    .X(_07106_));
 sky130_fd_sc_hd__or3_1 _13936_ (.A(_07104_),
    .B(_06971_),
    .C(_06930_),
    .X(_07107_));
 sky130_fd_sc_hd__a21bo_1 _13937_ (.A1(_07058_),
    .A2(_07106_),
    .B1_N(_07107_),
    .X(_07108_));
 sky130_fd_sc_hd__or2b_1 _13938_ (.A(_07088_),
    .B_N(_07096_),
    .X(_07109_));
 sky130_fd_sc_hd__a21bo_1 _13939_ (.A1(_06879_),
    .A2(_07097_),
    .B1_N(_07109_),
    .X(_07110_));
 sky130_fd_sc_hd__nand2_1 _13940_ (.A(_07065_),
    .B(_07085_),
    .Y(_07111_));
 sky130_fd_sc_hd__o21ai_1 _13941_ (.A1(_07086_),
    .A2(_07098_),
    .B1(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__or2b_1 _13942_ (.A(_07072_),
    .B_N(_07071_),
    .X(_07113_));
 sky130_fd_sc_hd__a21bo_1 _13943_ (.A1(_07073_),
    .A2(_07084_),
    .B1_N(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__nand2_1 _13944_ (.A(_06742_),
    .B(_06743_),
    .Y(_07115_));
 sky130_fd_sc_hd__nand2_1 _13945_ (.A(_07067_),
    .B(_07115_),
    .Y(_07116_));
 sky130_fd_sc_hd__or3_1 _13946_ (.A(_06942_),
    .B(_06718_),
    .C(_07116_),
    .X(_07117_));
 sky130_fd_sc_hd__o21ai_1 _13947_ (.A1(_06942_),
    .A2(_06718_),
    .B1(_07116_),
    .Y(_07118_));
 sky130_fd_sc_hd__and2_1 _13948_ (.A(_07117_),
    .B(_07118_),
    .X(_07119_));
 sky130_fd_sc_hd__a22o_1 _13949_ (.A1(_06741_),
    .A2(_07066_),
    .B1(_07069_),
    .B2(_07070_),
    .X(_07120_));
 sky130_fd_sc_hd__o22a_1 _13950_ (.A1(_06707_),
    .A2(_07078_),
    .B1(_06759_),
    .B2(_06722_),
    .X(_07121_));
 sky130_fd_sc_hd__xnor2_1 _13951_ (.A(_07120_),
    .B(_07121_),
    .Y(_07122_));
 sky130_fd_sc_hd__nand2_1 _13952_ (.A(_06721_),
    .B(_06708_),
    .Y(_07123_));
 sky130_fd_sc_hd__and2_1 _13953_ (.A(_06748_),
    .B(_06722_),
    .X(_07124_));
 sky130_fd_sc_hd__nor2_1 _13954_ (.A(_07123_),
    .B(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__xnor2_1 _13955_ (.A(_07122_),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__nand2_1 _13956_ (.A(_07119_),
    .B(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__or2_1 _13957_ (.A(_07119_),
    .B(_07126_),
    .X(_07128_));
 sky130_fd_sc_hd__and2_1 _13958_ (.A(_07127_),
    .B(_07128_),
    .X(_07129_));
 sky130_fd_sc_hd__xnor2_2 _13959_ (.A(_07114_),
    .B(_07129_),
    .Y(_07130_));
 sky130_fd_sc_hd__and2_1 _13960_ (.A(_07075_),
    .B(_07083_),
    .X(_07131_));
 sky130_fd_sc_hd__nor2_1 _13961_ (.A(_06732_),
    .B(_06769_),
    .Y(_07132_));
 sky130_fd_sc_hd__nand2_1 _13962_ (.A(_07090_),
    .B(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__nor2_1 _13963_ (.A(_06732_),
    .B(_06719_),
    .Y(_07134_));
 sky130_fd_sc_hd__inv_2 _13964_ (.A(_07134_),
    .Y(_07135_));
 sky130_fd_sc_hd__o21ai_1 _13965_ (.A1(_06687_),
    .A2(_06769_),
    .B1(_07135_),
    .Y(_07136_));
 sky130_fd_sc_hd__and2_1 _13966_ (.A(_07133_),
    .B(_07136_),
    .X(_07137_));
 sky130_fd_sc_hd__xnor2_1 _13967_ (.A(_07091_),
    .B(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__o21a_1 _13968_ (.A1(_07081_),
    .A2(_07131_),
    .B1(_07138_),
    .X(_07139_));
 sky130_fd_sc_hd__nor3_1 _13969_ (.A(_07081_),
    .B(_07131_),
    .C(_07138_),
    .Y(_07140_));
 sky130_fd_sc_hd__nor2_1 _13970_ (.A(_07139_),
    .B(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__xnor2_1 _13971_ (.A(_07094_),
    .B(_07141_),
    .Y(_07142_));
 sky130_fd_sc_hd__xor2_2 _13972_ (.A(_07130_),
    .B(_07142_),
    .X(_07143_));
 sky130_fd_sc_hd__xnor2_1 _13973_ (.A(_07112_),
    .B(_07143_),
    .Y(_07144_));
 sky130_fd_sc_hd__xor2_1 _13974_ (.A(_07110_),
    .B(_07144_),
    .X(_07145_));
 sky130_fd_sc_hd__and2b_1 _13975_ (.A_N(_07063_),
    .B(_07099_),
    .X(_07146_));
 sky130_fd_sc_hd__a21oi_1 _13976_ (.A1(_07060_),
    .A2(_07100_),
    .B1(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__xnor2_1 _13977_ (.A(_07145_),
    .B(_07147_),
    .Y(_07148_));
 sky130_fd_sc_hd__nor2_1 _13978_ (.A(_07101_),
    .B(_07103_),
    .Y(_07149_));
 sky130_fd_sc_hd__inv_2 _13979_ (.A(_07149_),
    .Y(_07150_));
 sky130_fd_sc_hd__or3_1 _13980_ (.A(_07104_),
    .B(_06888_),
    .C(_06927_),
    .X(_07151_));
 sky130_fd_sc_hd__nand2_1 _13981_ (.A(_07150_),
    .B(_07151_),
    .Y(_07152_));
 sky130_fd_sc_hd__xnor2_1 _13982_ (.A(_07148_),
    .B(_07152_),
    .Y(_07153_));
 sky130_fd_sc_hd__xnor2_1 _13983_ (.A(_07108_),
    .B(_07153_),
    .Y(_07154_));
 sky130_fd_sc_hd__xor2_1 _13984_ (.A(_07058_),
    .B(_07106_),
    .X(_07155_));
 sky130_fd_sc_hd__xnor2_1 _13985_ (.A(_07055_),
    .B(_07057_),
    .Y(_07156_));
 sky130_fd_sc_hd__and2b_1 _13986_ (.A_N(_07054_),
    .B(_07043_),
    .X(_07157_));
 sky130_fd_sc_hd__xnor2_2 _13987_ (.A(_07157_),
    .B(_07053_),
    .Y(_07158_));
 sky130_fd_sc_hd__nor2_1 _13988_ (.A(_07156_),
    .B(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__nor2_1 _13989_ (.A(_07155_),
    .B(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__nand2_1 _13990_ (.A(_07154_),
    .B(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__a2bb2o_1 _13991_ (.A1_N(_07148_),
    .A2_N(_07151_),
    .B1(_07153_),
    .B2(_07108_),
    .X(_07162_));
 sky130_fd_sc_hd__nor2_1 _13992_ (.A(_07145_),
    .B(_07147_),
    .Y(_07163_));
 sky130_fd_sc_hd__nor2_1 _13993_ (.A(_07150_),
    .B(_07148_),
    .Y(_07164_));
 sky130_fd_sc_hd__and2b_1 _13994_ (.A_N(_07144_),
    .B(_07110_),
    .X(_07165_));
 sky130_fd_sc_hd__a21oi_2 _13995_ (.A1(_07112_),
    .A2(_07143_),
    .B1(_07165_),
    .Y(_07166_));
 sky130_fd_sc_hd__nor2_1 _13996_ (.A(_07130_),
    .B(_07142_),
    .Y(_07167_));
 sky130_fd_sc_hd__a21o_1 _13997_ (.A1(_07114_),
    .A2(_07129_),
    .B1(_07167_),
    .X(_07168_));
 sky130_fd_sc_hd__nand2_1 _13998_ (.A(_06721_),
    .B(_06758_),
    .Y(_07169_));
 sky130_fd_sc_hd__o211a_1 _13999_ (.A1(_06718_),
    .A2(_06755_),
    .B1(_06738_),
    .C1(_06723_),
    .X(_07170_));
 sky130_fd_sc_hd__a211o_1 _14000_ (.A1(_06723_),
    .A2(_06738_),
    .B1(_06993_),
    .C1(_06718_),
    .X(_07171_));
 sky130_fd_sc_hd__and2b_1 _14001_ (.A_N(_07170_),
    .B(_07171_),
    .X(_07172_));
 sky130_fd_sc_hd__xnor2_1 _14002_ (.A(_07169_),
    .B(_07172_),
    .Y(_07173_));
 sky130_fd_sc_hd__or2_1 _14003_ (.A(_07117_),
    .B(_07173_),
    .X(_07174_));
 sky130_fd_sc_hd__nand2_1 _14004_ (.A(_07117_),
    .B(_07173_),
    .Y(_07175_));
 sky130_fd_sc_hd__nand2_1 _14005_ (.A(_07174_),
    .B(_07175_),
    .Y(_07176_));
 sky130_fd_sc_hd__xnor2_1 _14006_ (.A(_06710_),
    .B(_07176_),
    .Y(_07177_));
 sky130_fd_sc_hd__or3_1 _14007_ (.A(_06540_),
    .B(_06942_),
    .C(_07177_),
    .X(_07178_));
 sky130_fd_sc_hd__o21ai_1 _14008_ (.A1(_06540_),
    .A2(_06942_),
    .B1(_07177_),
    .Y(_07179_));
 sky130_fd_sc_hd__and2_1 _14009_ (.A(_07178_),
    .B(_07179_),
    .X(_07180_));
 sky130_fd_sc_hd__xor2_1 _14010_ (.A(_07127_),
    .B(_07180_),
    .X(_07181_));
 sky130_fd_sc_hd__and3_1 _14011_ (.A(_07089_),
    .B(_07090_),
    .C(_07137_),
    .X(_07182_));
 sky130_fd_sc_hd__nand2_1 _14012_ (.A(_07120_),
    .B(_07121_),
    .Y(_07183_));
 sky130_fd_sc_hd__o31a_1 _14013_ (.A1(_07123_),
    .A2(_07122_),
    .A3(_07124_),
    .B1(_07183_),
    .X(_07184_));
 sky130_fd_sc_hd__or2_1 _14014_ (.A(_06733_),
    .B(_06719_),
    .X(_07185_));
 sky130_fd_sc_hd__xor2_1 _14015_ (.A(_07132_),
    .B(_07185_),
    .X(_07186_));
 sky130_fd_sc_hd__nor2_1 _14016_ (.A(_07133_),
    .B(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__and2_1 _14017_ (.A(_07133_),
    .B(_07186_),
    .X(_07188_));
 sky130_fd_sc_hd__nor2_1 _14018_ (.A(_07187_),
    .B(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__xnor2_1 _14019_ (.A(_07184_),
    .B(_07189_),
    .Y(_07190_));
 sky130_fd_sc_hd__xnor2_1 _14020_ (.A(_07182_),
    .B(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__or2_1 _14021_ (.A(_07181_),
    .B(_07191_),
    .X(_07192_));
 sky130_fd_sc_hd__nand2_1 _14022_ (.A(_07181_),
    .B(_07191_),
    .Y(_07193_));
 sky130_fd_sc_hd__nand2_1 _14023_ (.A(_07192_),
    .B(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__xnor2_1 _14024_ (.A(_07168_),
    .B(_07194_),
    .Y(_07195_));
 sky130_fd_sc_hd__a21oi_1 _14025_ (.A1(_07094_),
    .A2(_07141_),
    .B1(_07139_),
    .Y(_07196_));
 sky130_fd_sc_hd__xnor2_2 _14026_ (.A(_07195_),
    .B(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__xnor2_2 _14027_ (.A(_07166_),
    .B(_07197_),
    .Y(_07198_));
 sky130_fd_sc_hd__or3_1 _14028_ (.A(_07163_),
    .B(_07164_),
    .C(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__o21ai_1 _14029_ (.A1(_07163_),
    .A2(_07164_),
    .B1(_07198_),
    .Y(_07200_));
 sky130_fd_sc_hd__and2_1 _14030_ (.A(_07199_),
    .B(_07200_),
    .X(_07201_));
 sky130_fd_sc_hd__xor2_2 _14031_ (.A(_07162_),
    .B(_07201_),
    .X(_07202_));
 sky130_fd_sc_hd__xnor2_1 _14032_ (.A(_07161_),
    .B(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__clkbuf_4 _14033_ (.A(_07203_),
    .X(_07204_));
 sky130_fd_sc_hd__or2_1 _14034_ (.A(_06720_),
    .B(_07204_),
    .X(_07205_));
 sky130_fd_sc_hd__buf_2 _14035_ (.A(_06769_),
    .X(_07206_));
 sky130_fd_sc_hd__or2_1 _14036_ (.A(_07154_),
    .B(_07160_),
    .X(_07207_));
 sky130_fd_sc_hd__nand2_1 _14037_ (.A(_07161_),
    .B(_07207_),
    .Y(_07208_));
 sky130_fd_sc_hd__clkbuf_4 _14038_ (.A(_07208_),
    .X(_07209_));
 sky130_fd_sc_hd__nor2_1 _14039_ (.A(_07206_),
    .B(_07209_),
    .Y(_07210_));
 sky130_fd_sc_hd__and2b_1 _14040_ (.A_N(_07205_),
    .B(_07210_),
    .X(_07211_));
 sky130_fd_sc_hd__or2_2 _14041_ (.A(_07161_),
    .B(_07202_),
    .X(_07212_));
 sky130_fd_sc_hd__a22o_2 _14042_ (.A1(_07164_),
    .A2(_07198_),
    .B1(_07201_),
    .B2(_07162_),
    .X(_07213_));
 sky130_fd_sc_hd__nand2_2 _14043_ (.A(_07163_),
    .B(_07198_),
    .Y(_07214_));
 sky130_fd_sc_hd__and2b_2 _14044_ (.A_N(_07166_),
    .B(_07197_),
    .X(_07215_));
 sky130_fd_sc_hd__and3_1 _14045_ (.A(_07168_),
    .B(_07192_),
    .C(_07193_),
    .X(_07216_));
 sky130_fd_sc_hd__and2b_1 _14046_ (.A_N(_07196_),
    .B(_07195_),
    .X(_07217_));
 sky130_fd_sc_hd__or2b_1 _14047_ (.A(_07127_),
    .B_N(_07180_),
    .X(_07218_));
 sky130_fd_sc_hd__nor2_1 _14048_ (.A(_06718_),
    .B(_06727_),
    .Y(_07219_));
 sky130_fd_sc_hd__nand2_1 _14049_ (.A(_06759_),
    .B(_07219_),
    .Y(_07220_));
 sky130_fd_sc_hd__or2_1 _14050_ (.A(_06759_),
    .B(_07219_),
    .X(_07221_));
 sky130_fd_sc_hd__nand2_1 _14051_ (.A(_07220_),
    .B(_07221_),
    .Y(_07222_));
 sky130_fd_sc_hd__xnor2_1 _14052_ (.A(_07178_),
    .B(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__o21a_1 _14053_ (.A1(_06710_),
    .A2(_07176_),
    .B1(_07174_),
    .X(_07224_));
 sky130_fd_sc_hd__or2_1 _14054_ (.A(_06733_),
    .B(_06769_),
    .X(_07225_));
 sky130_fd_sc_hd__nor3_1 _14055_ (.A(_06640_),
    .B(_06769_),
    .C(_07185_),
    .Y(_07226_));
 sky130_fd_sc_hd__or3_1 _14056_ (.A(_07135_),
    .B(_07225_),
    .C(_07226_),
    .X(_07227_));
 sky130_fd_sc_hd__o21a_1 _14057_ (.A1(_06640_),
    .A2(_06719_),
    .B1(_07225_),
    .X(_07228_));
 sky130_fd_sc_hd__o22ai_1 _14058_ (.A1(_07135_),
    .A2(_07225_),
    .B1(_07226_),
    .B2(_07228_),
    .Y(_07229_));
 sky130_fd_sc_hd__and2_1 _14059_ (.A(_07227_),
    .B(_07229_),
    .X(_07230_));
 sky130_fd_sc_hd__xnor2_1 _14060_ (.A(_07224_),
    .B(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__xnor2_1 _14061_ (.A(_07187_),
    .B(_07231_),
    .Y(_07232_));
 sky130_fd_sc_hd__or2_1 _14062_ (.A(_07223_),
    .B(_07232_),
    .X(_07233_));
 sky130_fd_sc_hd__nand2_1 _14063_ (.A(_07223_),
    .B(_07232_),
    .Y(_07234_));
 sky130_fd_sc_hd__nand2_1 _14064_ (.A(_07233_),
    .B(_07234_),
    .Y(_07235_));
 sky130_fd_sc_hd__a21oi_1 _14065_ (.A1(_07218_),
    .A2(_07192_),
    .B1(_07235_),
    .Y(_07236_));
 sky130_fd_sc_hd__and3_1 _14066_ (.A(_07218_),
    .B(_07192_),
    .C(_07235_),
    .X(_07237_));
 sky130_fd_sc_hd__or2_1 _14067_ (.A(_07236_),
    .B(_07237_),
    .X(_07238_));
 sky130_fd_sc_hd__or2b_1 _14068_ (.A(_07184_),
    .B_N(_07189_),
    .X(_07239_));
 sky130_fd_sc_hd__a21bo_1 _14069_ (.A1(_07182_),
    .A2(_07190_),
    .B1_N(_07239_),
    .X(_07240_));
 sky130_fd_sc_hd__xnor2_1 _14070_ (.A(_07238_),
    .B(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__o21a_2 _14071_ (.A1(_07216_),
    .A2(_07217_),
    .B1(_07241_),
    .X(_07242_));
 sky130_fd_sc_hd__nor3_1 _14072_ (.A(_07216_),
    .B(_07217_),
    .C(_07241_),
    .Y(_07243_));
 sky130_fd_sc_hd__nor2_2 _14073_ (.A(_07242_),
    .B(_07243_),
    .Y(_07244_));
 sky130_fd_sc_hd__xor2_4 _14074_ (.A(_07215_),
    .B(_07244_),
    .X(_07245_));
 sky130_fd_sc_hd__xnor2_4 _14075_ (.A(_07214_),
    .B(_07245_),
    .Y(_07246_));
 sky130_fd_sc_hd__xor2_4 _14076_ (.A(_07213_),
    .B(_07246_),
    .X(_07247_));
 sky130_fd_sc_hd__xnor2_4 _14077_ (.A(_07212_),
    .B(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__clkbuf_4 _14078_ (.A(_07248_),
    .X(_07249_));
 sky130_fd_sc_hd__o22ai_1 _14079_ (.A1(_06720_),
    .A2(_07249_),
    .B1(_07204_),
    .B2(_07206_),
    .Y(_07250_));
 sky130_fd_sc_hd__o31a_1 _14080_ (.A1(_07206_),
    .A2(_07249_),
    .A3(_07205_),
    .B1(_07250_),
    .X(_07251_));
 sky130_fd_sc_hd__clkbuf_4 _14081_ (.A(_06942_),
    .X(_07252_));
 sky130_fd_sc_hd__clkbuf_4 _14082_ (.A(_06857_),
    .X(_07253_));
 sky130_fd_sc_hd__or2_2 _14083_ (.A(_07212_),
    .B(_07247_),
    .X(_07254_));
 sky130_fd_sc_hd__and3_1 _14084_ (.A(_07163_),
    .B(_07198_),
    .C(_07245_),
    .X(_07255_));
 sky130_fd_sc_hd__a21oi_2 _14085_ (.A1(_07213_),
    .A2(_07246_),
    .B1(_07255_),
    .Y(_07256_));
 sky130_fd_sc_hd__nand2_1 _14086_ (.A(_07215_),
    .B(_07244_),
    .Y(_07257_));
 sky130_fd_sc_hd__and2b_1 _14087_ (.A_N(_07238_),
    .B(_07240_),
    .X(_07258_));
 sky130_fd_sc_hd__o21ai_1 _14088_ (.A1(_07178_),
    .A2(_07222_),
    .B1(_07233_),
    .Y(_07259_));
 sky130_fd_sc_hd__nor2_1 _14089_ (.A(_06722_),
    .B(_07123_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand2_1 _14090_ (.A(_07260_),
    .B(_07221_),
    .Y(_07261_));
 sky130_fd_sc_hd__o22a_1 _14091_ (.A1(_06718_),
    .A2(_07078_),
    .B1(_06727_),
    .B2(_06540_),
    .X(_07262_));
 sky130_fd_sc_hd__a31o_1 _14092_ (.A1(_07067_),
    .A2(_06758_),
    .A3(_07219_),
    .B1(_07262_),
    .X(_07263_));
 sky130_fd_sc_hd__a21o_1 _14093_ (.A1(_07220_),
    .A2(_07261_),
    .B1(_07263_),
    .X(_07264_));
 sky130_fd_sc_hd__nand3_1 _14094_ (.A(_07220_),
    .B(_07261_),
    .C(_07263_),
    .Y(_07265_));
 sky130_fd_sc_hd__nand2_1 _14095_ (.A(_07264_),
    .B(_07265_),
    .Y(_07266_));
 sky130_fd_sc_hd__o22a_1 _14096_ (.A1(_06640_),
    .A2(_06769_),
    .B1(_06720_),
    .B2(_06722_),
    .X(_07267_));
 sky130_fd_sc_hd__or4_1 _14097_ (.A(_06722_),
    .B(_06640_),
    .C(_06769_),
    .D(_06720_),
    .X(_07268_));
 sky130_fd_sc_hd__and2_1 _14098_ (.A(_07260_),
    .B(_07222_),
    .X(_07269_));
 sky130_fd_sc_hd__inv_2 _14099_ (.A(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__or4bb_1 _14100_ (.A(_07226_),
    .B(_07267_),
    .C_N(_07268_),
    .D_N(_07270_),
    .X(_07271_));
 sky130_fd_sc_hd__xnor2_1 _14101_ (.A(_07227_),
    .B(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__or2_1 _14102_ (.A(_07266_),
    .B(_07272_),
    .X(_07273_));
 sky130_fd_sc_hd__nand2_1 _14103_ (.A(_07266_),
    .B(_07272_),
    .Y(_07274_));
 sky130_fd_sc_hd__and2_1 _14104_ (.A(_07273_),
    .B(_07274_),
    .X(_07275_));
 sky130_fd_sc_hd__xnor2_1 _14105_ (.A(_07259_),
    .B(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__or2b_1 _14106_ (.A(_07224_),
    .B_N(_07230_),
    .X(_07277_));
 sky130_fd_sc_hd__a21bo_1 _14107_ (.A1(_07187_),
    .A2(_07231_),
    .B1_N(_07277_),
    .X(_07278_));
 sky130_fd_sc_hd__xnor2_1 _14108_ (.A(_07276_),
    .B(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__o21ai_1 _14109_ (.A1(_07236_),
    .A2(_07258_),
    .B1(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__or3_1 _14110_ (.A(_07236_),
    .B(_07258_),
    .C(_07279_),
    .X(_07281_));
 sky130_fd_sc_hd__and2_1 _14111_ (.A(_07280_),
    .B(_07281_),
    .X(_07282_));
 sky130_fd_sc_hd__xor2_4 _14112_ (.A(_07242_),
    .B(_07282_),
    .X(_07283_));
 sky130_fd_sc_hd__xnor2_2 _14113_ (.A(_07257_),
    .B(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__xnor2_4 _14114_ (.A(_07256_),
    .B(_07284_),
    .Y(_07285_));
 sky130_fd_sc_hd__and2_1 _14115_ (.A(_07213_),
    .B(_07246_),
    .X(_07286_));
 sky130_fd_sc_hd__and2b_1 _14116_ (.A_N(_07276_),
    .B(_07278_),
    .X(_07287_));
 sky130_fd_sc_hd__a21oi_1 _14117_ (.A1(_07259_),
    .A2(_07275_),
    .B1(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__or3_1 _14118_ (.A(_06540_),
    .B(_07078_),
    .C(_07219_),
    .X(_07289_));
 sky130_fd_sc_hd__and2_1 _14119_ (.A(_06723_),
    .B(_07268_),
    .X(_07290_));
 sky130_fd_sc_hd__xnor2_1 _14120_ (.A(_07264_),
    .B(_07290_),
    .Y(_07291_));
 sky130_fd_sc_hd__nor2_1 _14121_ (.A(_07226_),
    .B(_07291_),
    .Y(_07292_));
 sky130_fd_sc_hd__xnor2_1 _14122_ (.A(_07289_),
    .B(_07292_),
    .Y(_07293_));
 sky130_fd_sc_hd__o211a_1 _14123_ (.A1(_07227_),
    .A2(_07271_),
    .B1(_07273_),
    .C1(_07270_),
    .X(_07294_));
 sky130_fd_sc_hd__xnor2_1 _14124_ (.A(_07293_),
    .B(_07294_),
    .Y(_07295_));
 sky130_fd_sc_hd__xnor2_1 _14125_ (.A(_07288_),
    .B(_07295_),
    .Y(_07296_));
 sky130_fd_sc_hd__nor2_1 _14126_ (.A(_07280_),
    .B(_07296_),
    .Y(_07297_));
 sky130_fd_sc_hd__a221o_1 _14127_ (.A1(_07242_),
    .A2(_07282_),
    .B1(_07296_),
    .B2(_07280_),
    .C1(_07297_),
    .X(_07298_));
 sky130_fd_sc_hd__inv_2 _14128_ (.A(_07257_),
    .Y(_07299_));
 sky130_fd_sc_hd__o21a_1 _14129_ (.A1(_07299_),
    .A2(_07255_),
    .B1(_07283_),
    .X(_07300_));
 sky130_fd_sc_hd__a211o_1 _14130_ (.A1(_07286_),
    .A2(_07284_),
    .B1(_07298_),
    .C1(_07300_),
    .X(_07301_));
 sky130_fd_sc_hd__o21ai_2 _14131_ (.A1(_07254_),
    .A2(_07285_),
    .B1(_07301_),
    .Y(_07302_));
 sky130_fd_sc_hd__clkbuf_2 _14132_ (.A(_07302_),
    .X(_07303_));
 sky130_fd_sc_hd__or3_1 _14133_ (.A(_07252_),
    .B(_07253_),
    .C(_07303_),
    .X(_07304_));
 sky130_fd_sc_hd__or2_2 _14134_ (.A(_06993_),
    .B(_07303_),
    .X(_07305_));
 sky130_fd_sc_hd__buf_2 _14135_ (.A(_06727_),
    .X(_07306_));
 sky130_fd_sc_hd__nor2_1 _14136_ (.A(_07306_),
    .B(_07303_),
    .Y(_07307_));
 sky130_fd_sc_hd__xnor2_1 _14137_ (.A(_07305_),
    .B(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__xor2_4 _14138_ (.A(_07254_),
    .B(_07285_),
    .X(_07309_));
 sky130_fd_sc_hd__buf_2 _14139_ (.A(_07309_),
    .X(_07310_));
 sky130_fd_sc_hd__and2_1 _14140_ (.A(_06758_),
    .B(_07310_),
    .X(_07311_));
 sky130_fd_sc_hd__xor2_1 _14141_ (.A(_07308_),
    .B(_07311_),
    .X(_07312_));
 sky130_fd_sc_hd__or2b_1 _14142_ (.A(_07304_),
    .B_N(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__xor2_1 _14143_ (.A(_07304_),
    .B(_07312_),
    .X(_07314_));
 sky130_fd_sc_hd__nand2_1 _14144_ (.A(_06738_),
    .B(_07310_),
    .Y(_07315_));
 sky130_fd_sc_hd__buf_2 _14145_ (.A(_07078_),
    .X(_07316_));
 sky130_fd_sc_hd__xor2_1 _14146_ (.A(_07305_),
    .B(_07315_),
    .X(_07317_));
 sky130_fd_sc_hd__or3b_1 _14147_ (.A(_07316_),
    .B(_07249_),
    .C_N(_07317_),
    .X(_07318_));
 sky130_fd_sc_hd__o21a_1 _14148_ (.A1(_07305_),
    .A2(_07315_),
    .B1(_07318_),
    .X(_07319_));
 sky130_fd_sc_hd__or2_1 _14149_ (.A(_07314_),
    .B(_07319_),
    .X(_07320_));
 sky130_fd_sc_hd__nand2_1 _14150_ (.A(_06775_),
    .B(_07310_),
    .Y(_07321_));
 sky130_fd_sc_hd__or3b_1 _14151_ (.A(_07206_),
    .B(_07249_),
    .C_N(_07205_),
    .X(_07322_));
 sky130_fd_sc_hd__xnor2_1 _14152_ (.A(_07321_),
    .B(_07322_),
    .Y(_07323_));
 sky130_fd_sc_hd__a21oi_1 _14153_ (.A1(_07313_),
    .A2(_07320_),
    .B1(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__and3_1 _14154_ (.A(_07313_),
    .B(_07320_),
    .C(_07323_),
    .X(_07325_));
 sky130_fd_sc_hd__nor2_1 _14155_ (.A(_07324_),
    .B(_07325_),
    .Y(_07326_));
 sky130_fd_sc_hd__a31o_1 _14156_ (.A1(_07211_),
    .A2(_07251_),
    .A3(_07326_),
    .B1(_07324_),
    .X(_07327_));
 sky130_fd_sc_hd__or2_1 _14157_ (.A(_07306_),
    .B(_07305_),
    .X(_07328_));
 sky130_fd_sc_hd__nor2_1 _14158_ (.A(_07316_),
    .B(_07303_),
    .Y(_07329_));
 sky130_fd_sc_hd__nand2_1 _14159_ (.A(_07308_),
    .B(_07329_),
    .Y(_07330_));
 sky130_fd_sc_hd__buf_2 _14160_ (.A(_07303_),
    .X(_07331_));
 sky130_fd_sc_hd__or3_1 _14161_ (.A(_07316_),
    .B(_07306_),
    .C(_07331_),
    .X(_07332_));
 sky130_fd_sc_hd__a21bo_1 _14162_ (.A1(_07328_),
    .A2(_07330_),
    .B1_N(_07332_),
    .X(_07333_));
 sky130_fd_sc_hd__a311o_1 _14163_ (.A1(_07067_),
    .A2(_06759_),
    .A3(_07331_),
    .B1(_07307_),
    .C1(_07329_),
    .X(_07334_));
 sky130_fd_sc_hd__a21oi_1 _14164_ (.A1(_07333_),
    .A2(_07334_),
    .B1(_06540_),
    .Y(_07335_));
 sky130_fd_sc_hd__or2b_1 _14165_ (.A(_07264_),
    .B_N(_07290_),
    .X(_07336_));
 sky130_fd_sc_hd__nor2_1 _14166_ (.A(_06720_),
    .B(_07331_),
    .Y(_07337_));
 sky130_fd_sc_hd__or2b_1 _14167_ (.A(_07206_),
    .B_N(_07310_),
    .X(_07338_));
 sky130_fd_sc_hd__a21o_1 _14168_ (.A1(_07249_),
    .A2(_07337_),
    .B1(_07338_),
    .X(_07339_));
 sky130_fd_sc_hd__nand2_1 _14169_ (.A(_07336_),
    .B(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__xor2_1 _14170_ (.A(_07335_),
    .B(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__nand2_1 _14171_ (.A(_07211_),
    .B(_07251_),
    .Y(_07342_));
 sky130_fd_sc_hd__xnor2_1 _14172_ (.A(_07342_),
    .B(_07326_),
    .Y(_07343_));
 sky130_fd_sc_hd__nor2_1 _14173_ (.A(_07252_),
    .B(_07303_),
    .Y(_07344_));
 sky130_fd_sc_hd__a21o_1 _14174_ (.A1(_07115_),
    .A2(_07331_),
    .B1(_07344_),
    .X(_07345_));
 sky130_fd_sc_hd__xor2_1 _14175_ (.A(_07314_),
    .B(_07319_),
    .X(_07346_));
 sky130_fd_sc_hd__nand2_1 _14176_ (.A(_07345_),
    .B(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__or2_1 _14177_ (.A(_07308_),
    .B(_07329_),
    .X(_07348_));
 sky130_fd_sc_hd__o21ai_1 _14178_ (.A1(_07311_),
    .A2(_07330_),
    .B1(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__nand2_1 _14179_ (.A(_07328_),
    .B(_07349_),
    .Y(_07350_));
 sky130_fd_sc_hd__a22oi_2 _14180_ (.A1(_06854_),
    .A2(_07331_),
    .B1(_07350_),
    .B2(_07336_),
    .Y(_07351_));
 sky130_fd_sc_hd__nor2_1 _14181_ (.A(_07347_),
    .B(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__and2_1 _14182_ (.A(_07347_),
    .B(_07351_),
    .X(_07353_));
 sky130_fd_sc_hd__nor2_1 _14183_ (.A(_07352_),
    .B(_07353_),
    .Y(_07354_));
 sky130_fd_sc_hd__a21oi_1 _14184_ (.A1(_07343_),
    .A2(_07354_),
    .B1(_07352_),
    .Y(_07355_));
 sky130_fd_sc_hd__xor2_1 _14185_ (.A(_07341_),
    .B(_07355_),
    .X(_07356_));
 sky130_fd_sc_hd__xnor2_1 _14186_ (.A(_07327_),
    .B(_07356_),
    .Y(_07357_));
 sky130_fd_sc_hd__xnor2_1 _14187_ (.A(_07343_),
    .B(_07354_),
    .Y(_07358_));
 sky130_fd_sc_hd__and2_1 _14188_ (.A(_07155_),
    .B(_07159_),
    .X(_07359_));
 sky130_fd_sc_hd__or2_1 _14189_ (.A(_07160_),
    .B(_07359_),
    .X(_07360_));
 sky130_fd_sc_hd__clkbuf_4 _14190_ (.A(_07360_),
    .X(_07361_));
 sky130_fd_sc_hd__nor2_1 _14191_ (.A(_06720_),
    .B(_07361_),
    .Y(_07362_));
 sky130_fd_sc_hd__and3_1 _14192_ (.A(_07205_),
    .B(_07210_),
    .C(_07362_),
    .X(_07363_));
 sky130_fd_sc_hd__or2_1 _14193_ (.A(_07211_),
    .B(_07251_),
    .X(_07364_));
 sky130_fd_sc_hd__nand2_1 _14194_ (.A(_07342_),
    .B(_07364_),
    .Y(_07365_));
 sky130_fd_sc_hd__clkbuf_2 _14195_ (.A(_07302_),
    .X(_07366_));
 sky130_fd_sc_hd__or3_2 _14196_ (.A(_07253_),
    .B(_07045_),
    .C(_07366_),
    .X(_07367_));
 sky130_fd_sc_hd__a21oi_1 _14197_ (.A1(_07253_),
    .A2(_07045_),
    .B1(_07366_),
    .Y(_07368_));
 sky130_fd_sc_hd__and2_1 _14198_ (.A(_07367_),
    .B(_07368_),
    .X(_07369_));
 sky130_fd_sc_hd__nand2_1 _14199_ (.A(_07344_),
    .B(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__nand2_1 _14200_ (.A(_07367_),
    .B(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__o21bai_1 _14201_ (.A1(_07316_),
    .A2(_07249_),
    .B1_N(_07317_),
    .Y(_07372_));
 sky130_fd_sc_hd__nand2_1 _14202_ (.A(_07318_),
    .B(_07372_),
    .Y(_07373_));
 sky130_fd_sc_hd__xnor2_1 _14203_ (.A(_07371_),
    .B(_07373_),
    .Y(_07374_));
 sky130_fd_sc_hd__or2_1 _14204_ (.A(_07316_),
    .B(_07204_),
    .X(_07375_));
 sky130_fd_sc_hd__o2bb2a_1 _14205_ (.A1_N(_06759_),
    .A2_N(_07310_),
    .B1(_07249_),
    .B2(_07306_),
    .X(_07376_));
 sky130_fd_sc_hd__nor2_1 _14206_ (.A(_07375_),
    .B(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__a32o_1 _14207_ (.A1(_07318_),
    .A2(_07371_),
    .A3(_07372_),
    .B1(_07374_),
    .B2(_07377_),
    .X(_07378_));
 sky130_fd_sc_hd__xnor2_1 _14208_ (.A(_07365_),
    .B(_07378_),
    .Y(_07379_));
 sky130_fd_sc_hd__xor2_1 _14209_ (.A(_07363_),
    .B(_07379_),
    .X(_07380_));
 sky130_fd_sc_hd__nor2_1 _14210_ (.A(_07253_),
    .B(_07331_),
    .Y(_07381_));
 sky130_fd_sc_hd__a311o_1 _14211_ (.A1(_07067_),
    .A2(_06741_),
    .A3(_07331_),
    .B1(_07344_),
    .C1(_07381_),
    .X(_07382_));
 sky130_fd_sc_hd__and2_1 _14212_ (.A(_07304_),
    .B(_07382_),
    .X(_07383_));
 sky130_fd_sc_hd__xor2_2 _14213_ (.A(_07377_),
    .B(_07374_),
    .X(_07384_));
 sky130_fd_sc_hd__nand2_1 _14214_ (.A(_07383_),
    .B(_07384_),
    .Y(_07385_));
 sky130_fd_sc_hd__or2_1 _14215_ (.A(_07345_),
    .B(_07346_),
    .X(_07386_));
 sky130_fd_sc_hd__and2_1 _14216_ (.A(_07347_),
    .B(_07386_),
    .X(_07387_));
 sky130_fd_sc_hd__xnor2_1 _14217_ (.A(_07385_),
    .B(_07387_),
    .Y(_07388_));
 sky130_fd_sc_hd__and3_1 _14218_ (.A(_07383_),
    .B(_07384_),
    .C(_07387_),
    .X(_07389_));
 sky130_fd_sc_hd__a21oi_1 _14219_ (.A1(_07380_),
    .A2(_07388_),
    .B1(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__xnor2_1 _14220_ (.A(_07358_),
    .B(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__a32o_1 _14221_ (.A1(_07342_),
    .A2(_07364_),
    .A3(_07378_),
    .B1(_07379_),
    .B2(_07363_),
    .X(_07392_));
 sky130_fd_sc_hd__or2b_1 _14222_ (.A(_07391_),
    .B_N(_07392_),
    .X(_07393_));
 sky130_fd_sc_hd__o21a_1 _14223_ (.A1(_07358_),
    .A2(_07390_),
    .B1(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__nor2_1 _14224_ (.A(_07357_),
    .B(_07394_),
    .Y(_07395_));
 sky130_fd_sc_hd__and2_1 _14225_ (.A(_07338_),
    .B(_07337_),
    .X(_07396_));
 sky130_fd_sc_hd__or3b_1 _14226_ (.A(_07331_),
    .B(_07396_),
    .C_N(_07333_),
    .X(_07397_));
 sky130_fd_sc_hd__nand2_2 _14227_ (.A(_07067_),
    .B(_07366_),
    .Y(_07398_));
 sky130_fd_sc_hd__nor2_1 _14228_ (.A(_07306_),
    .B(_07398_),
    .Y(_07399_));
 sky130_fd_sc_hd__o21ai_1 _14229_ (.A1(_07329_),
    .A2(_07399_),
    .B1(_07332_),
    .Y(_07400_));
 sky130_fd_sc_hd__or2_1 _14230_ (.A(_07397_),
    .B(_07400_),
    .X(_07401_));
 sky130_fd_sc_hd__nand3b_2 _14231_ (.A_N(_07335_),
    .B(_07340_),
    .C(_07401_),
    .Y(_07402_));
 sky130_fd_sc_hd__nand2_1 _14232_ (.A(_07397_),
    .B(_07400_),
    .Y(_07403_));
 sky130_fd_sc_hd__a21oi_1 _14233_ (.A1(_07402_),
    .A2(_07403_),
    .B1(_07396_),
    .Y(_07404_));
 sky130_fd_sc_hd__nor2_1 _14234_ (.A(_07341_),
    .B(_07355_),
    .Y(_07405_));
 sky130_fd_sc_hd__a21oi_1 _14235_ (.A1(_07327_),
    .A2(_07356_),
    .B1(_07405_),
    .Y(_07406_));
 sky130_fd_sc_hd__or2_1 _14236_ (.A(_07404_),
    .B(_07406_),
    .X(_07407_));
 sky130_fd_sc_hd__nand2_1 _14237_ (.A(_07404_),
    .B(_07406_),
    .Y(_07408_));
 sky130_fd_sc_hd__and3_1 _14238_ (.A(_07395_),
    .B(_07407_),
    .C(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__and2_1 _14239_ (.A(_07407_),
    .B(_07408_),
    .X(_07410_));
 sky130_fd_sc_hd__nor2_1 _14240_ (.A(_07395_),
    .B(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__nor2_1 _14241_ (.A(_07409_),
    .B(_07411_),
    .Y(_07412_));
 sky130_fd_sc_hd__xor2_2 _14242_ (.A(_07392_),
    .B(_07391_),
    .X(_07413_));
 sky130_fd_sc_hd__xnor2_1 _14243_ (.A(_07380_),
    .B(_07388_),
    .Y(_07414_));
 sky130_fd_sc_hd__xnor2_1 _14244_ (.A(_07383_),
    .B(_07384_),
    .Y(_07415_));
 sky130_fd_sc_hd__or2_1 _14245_ (.A(_07344_),
    .B(_07369_),
    .X(_07416_));
 sky130_fd_sc_hd__clkbuf_4 _14246_ (.A(_06785_),
    .X(_07417_));
 sky130_fd_sc_hd__nor2_1 _14247_ (.A(_07417_),
    .B(_07398_),
    .Y(_07418_));
 sky130_fd_sc_hd__a211o_1 _14248_ (.A1(_07370_),
    .A2(_07416_),
    .B1(_07418_),
    .C1(_06540_),
    .X(_07419_));
 sky130_fd_sc_hd__and2_1 _14249_ (.A(_06854_),
    .B(_07309_),
    .X(_07420_));
 sky130_fd_sc_hd__nand3_1 _14250_ (.A(_07367_),
    .B(_07368_),
    .C(_07420_),
    .Y(_07421_));
 sky130_fd_sc_hd__a21o_1 _14251_ (.A1(_07367_),
    .A2(_07368_),
    .B1(_07420_),
    .X(_07422_));
 sky130_fd_sc_hd__clkbuf_4 _14252_ (.A(_06792_),
    .X(_07423_));
 sky130_fd_sc_hd__or2_1 _14253_ (.A(_07417_),
    .B(_07366_),
    .X(_07424_));
 sky130_fd_sc_hd__o21ai_1 _14254_ (.A1(_07423_),
    .A2(_07398_),
    .B1(_07424_),
    .Y(_07425_));
 sky130_fd_sc_hd__and3b_1 _14255_ (.A_N(_07303_),
    .B(_06807_),
    .C(_06808_),
    .X(_07426_));
 sky130_fd_sc_hd__a31o_1 _14256_ (.A1(_07421_),
    .A2(_07422_),
    .A3(_07425_),
    .B1(_07426_),
    .X(_07427_));
 sky130_fd_sc_hd__xnor2_1 _14257_ (.A(_07375_),
    .B(_07376_),
    .Y(_07428_));
 sky130_fd_sc_hd__a21o_1 _14258_ (.A1(_07367_),
    .A2(_07421_),
    .B1(_07428_),
    .X(_07429_));
 sky130_fd_sc_hd__nand3_1 _14259_ (.A(_07367_),
    .B(_07421_),
    .C(_07428_),
    .Y(_07430_));
 sky130_fd_sc_hd__nand2_1 _14260_ (.A(_07429_),
    .B(_07430_),
    .Y(_07431_));
 sky130_fd_sc_hd__or2_2 _14261_ (.A(_07306_),
    .B(_07203_),
    .X(_07432_));
 sky130_fd_sc_hd__or2_1 _14262_ (.A(_07316_),
    .B(_07209_),
    .X(_07433_));
 sky130_fd_sc_hd__nor2_1 _14263_ (.A(_06993_),
    .B(_07248_),
    .Y(_07434_));
 sky130_fd_sc_hd__xnor2_1 _14264_ (.A(_07432_),
    .B(_07434_),
    .Y(_07435_));
 sky130_fd_sc_hd__or2b_1 _14265_ (.A(_07433_),
    .B_N(_07435_),
    .X(_07436_));
 sky130_fd_sc_hd__o31a_1 _14266_ (.A1(_06993_),
    .A2(_07249_),
    .A3(_07432_),
    .B1(_07436_),
    .X(_07437_));
 sky130_fd_sc_hd__xor2_1 _14267_ (.A(_07431_),
    .B(_07437_),
    .X(_07438_));
 sky130_fd_sc_hd__xor2_1 _14268_ (.A(_07419_),
    .B(_07427_),
    .X(_07439_));
 sky130_fd_sc_hd__and2_1 _14269_ (.A(_07438_),
    .B(_07439_),
    .X(_07440_));
 sky130_fd_sc_hd__a21oi_1 _14270_ (.A1(_07419_),
    .A2(_07427_),
    .B1(_07440_),
    .Y(_07441_));
 sky130_fd_sc_hd__and2_1 _14271_ (.A(_07156_),
    .B(_07158_),
    .X(_07442_));
 sky130_fd_sc_hd__nor2_1 _14272_ (.A(_07159_),
    .B(_07442_),
    .Y(_07443_));
 sky130_fd_sc_hd__clkbuf_4 _14273_ (.A(_07443_),
    .X(_07444_));
 sky130_fd_sc_hd__nor2_1 _14274_ (.A(_07206_),
    .B(_07444_),
    .Y(_07445_));
 sky130_fd_sc_hd__nand2_1 _14275_ (.A(_07362_),
    .B(_07445_),
    .Y(_07446_));
 sky130_fd_sc_hd__nand2_1 _14276_ (.A(_07210_),
    .B(_07362_),
    .Y(_07447_));
 sky130_fd_sc_hd__nor2_1 _14277_ (.A(_06720_),
    .B(_07209_),
    .Y(_07448_));
 sky130_fd_sc_hd__nor2_1 _14278_ (.A(_07206_),
    .B(_07361_),
    .Y(_07449_));
 sky130_fd_sc_hd__or2_1 _14279_ (.A(_07448_),
    .B(_07449_),
    .X(_07450_));
 sky130_fd_sc_hd__a21oi_1 _14280_ (.A1(_07447_),
    .A2(_07450_),
    .B1(_06540_),
    .Y(_07451_));
 sky130_fd_sc_hd__or2_1 _14281_ (.A(_07446_),
    .B(_07451_),
    .X(_07452_));
 sky130_fd_sc_hd__o21a_1 _14282_ (.A1(_07206_),
    .A2(_07209_),
    .B1(_07205_),
    .X(_07453_));
 sky130_fd_sc_hd__o2bb2a_1 _14283_ (.A1_N(_07448_),
    .A2_N(_07449_),
    .B1(_07453_),
    .B2(_07211_),
    .X(_07454_));
 sky130_fd_sc_hd__or2_1 _14284_ (.A(_07363_),
    .B(_07454_),
    .X(_07455_));
 sky130_fd_sc_hd__o21a_1 _14285_ (.A1(_07431_),
    .A2(_07437_),
    .B1(_07429_),
    .X(_07456_));
 sky130_fd_sc_hd__xor2_1 _14286_ (.A(_07455_),
    .B(_07456_),
    .X(_07457_));
 sky130_fd_sc_hd__xnor2_1 _14287_ (.A(_07452_),
    .B(_07457_),
    .Y(_07458_));
 sky130_fd_sc_hd__xor2_1 _14288_ (.A(_07415_),
    .B(_07441_),
    .X(_07459_));
 sky130_fd_sc_hd__nand2_1 _14289_ (.A(_07458_),
    .B(_07459_),
    .Y(_07460_));
 sky130_fd_sc_hd__o21a_1 _14290_ (.A1(_07415_),
    .A2(_07441_),
    .B1(_07460_),
    .X(_07461_));
 sky130_fd_sc_hd__xnor2_1 _14291_ (.A(_07414_),
    .B(_07461_),
    .Y(_07462_));
 sky130_fd_sc_hd__or2b_1 _14292_ (.A(_07452_),
    .B_N(_07457_),
    .X(_07463_));
 sky130_fd_sc_hd__o21ai_2 _14293_ (.A1(_07455_),
    .A2(_07456_),
    .B1(_07463_),
    .Y(_07464_));
 sky130_fd_sc_hd__or2b_1 _14294_ (.A(_07462_),
    .B_N(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__o21a_1 _14295_ (.A1(_07414_),
    .A2(_07461_),
    .B1(_07465_),
    .X(_07466_));
 sky130_fd_sc_hd__nor2_1 _14296_ (.A(_07413_),
    .B(_07466_),
    .Y(_07467_));
 sky130_fd_sc_hd__and2_1 _14297_ (.A(_07357_),
    .B(_07394_),
    .X(_07468_));
 sky130_fd_sc_hd__nor2_1 _14298_ (.A(_07395_),
    .B(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__and2_1 _14299_ (.A(_07467_),
    .B(_07469_),
    .X(_07470_));
 sky130_fd_sc_hd__xor2_1 _14300_ (.A(_07412_),
    .B(_07470_),
    .X(_07471_));
 sky130_fd_sc_hd__xor2_1 _14301_ (.A(_07467_),
    .B(_07469_),
    .X(_07472_));
 sky130_fd_sc_hd__xor2_2 _14302_ (.A(_07464_),
    .B(_07462_),
    .X(_07473_));
 sky130_fd_sc_hd__or2_1 _14303_ (.A(_07458_),
    .B(_07459_),
    .X(_07474_));
 sky130_fd_sc_hd__nand2_1 _14304_ (.A(_07460_),
    .B(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__clkbuf_4 _14305_ (.A(_07158_),
    .X(_07476_));
 sky130_fd_sc_hd__nor2_1 _14306_ (.A(_06720_),
    .B(_07476_),
    .Y(_07477_));
 sky130_fd_sc_hd__and2_1 _14307_ (.A(_07445_),
    .B(_07477_),
    .X(_07478_));
 sky130_fd_sc_hd__nand2_1 _14308_ (.A(_07446_),
    .B(_07478_),
    .Y(_07479_));
 sky130_fd_sc_hd__nand2_1 _14309_ (.A(_07446_),
    .B(_07451_),
    .Y(_07480_));
 sky130_fd_sc_hd__nand2_1 _14310_ (.A(_07452_),
    .B(_07480_),
    .Y(_07481_));
 sky130_fd_sc_hd__nor2_1 _14311_ (.A(_07045_),
    .B(_07366_),
    .Y(_07482_));
 sky130_fd_sc_hd__and2_1 _14312_ (.A(_07115_),
    .B(_07309_),
    .X(_07483_));
 sky130_fd_sc_hd__xnor2_1 _14313_ (.A(_07482_),
    .B(_07483_),
    .Y(_07484_));
 sky130_fd_sc_hd__nand2_1 _14314_ (.A(_07482_),
    .B(_07483_),
    .Y(_07485_));
 sky130_fd_sc_hd__o31ai_2 _14315_ (.A1(_07252_),
    .A2(_07249_),
    .A3(_07484_),
    .B1(_07485_),
    .Y(_07486_));
 sky130_fd_sc_hd__xnor2_1 _14316_ (.A(_07433_),
    .B(_07435_),
    .Y(_07487_));
 sky130_fd_sc_hd__xnor2_1 _14317_ (.A(_07486_),
    .B(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__or2_1 _14318_ (.A(_06993_),
    .B(_07208_),
    .X(_07489_));
 sky130_fd_sc_hd__or2_1 _14319_ (.A(_07316_),
    .B(_07360_),
    .X(_07490_));
 sky130_fd_sc_hd__nor2_1 _14320_ (.A(_07306_),
    .B(_07208_),
    .Y(_07491_));
 sky130_fd_sc_hd__o21bai_1 _14321_ (.A1(_06993_),
    .A2(_07204_),
    .B1_N(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__o21ai_1 _14322_ (.A1(_07432_),
    .A2(_07489_),
    .B1(_07492_),
    .Y(_07493_));
 sky130_fd_sc_hd__o22a_1 _14323_ (.A1(_07432_),
    .A2(_07489_),
    .B1(_07490_),
    .B2(_07493_),
    .X(_07494_));
 sky130_fd_sc_hd__nand2_1 _14324_ (.A(_07486_),
    .B(_07487_),
    .Y(_07495_));
 sky130_fd_sc_hd__o21a_1 _14325_ (.A1(_07488_),
    .A2(_07494_),
    .B1(_07495_),
    .X(_07496_));
 sky130_fd_sc_hd__xor2_1 _14326_ (.A(_07481_),
    .B(_07496_),
    .X(_07497_));
 sky130_fd_sc_hd__xnor2_1 _14327_ (.A(_07479_),
    .B(_07497_),
    .Y(_07498_));
 sky130_fd_sc_hd__xnor2_1 _14328_ (.A(_07438_),
    .B(_07439_),
    .Y(_07499_));
 sky130_fd_sc_hd__xor2_1 _14329_ (.A(_07488_),
    .B(_07494_),
    .X(_07500_));
 sky130_fd_sc_hd__nand2_1 _14330_ (.A(_07421_),
    .B(_07422_),
    .Y(_07501_));
 sky130_fd_sc_hd__or2b_1 _14331_ (.A(_07426_),
    .B_N(_07425_),
    .X(_07502_));
 sky130_fd_sc_hd__xnor2_1 _14332_ (.A(_07501_),
    .B(_07502_),
    .Y(_07503_));
 sky130_fd_sc_hd__nor2_1 _14333_ (.A(_07252_),
    .B(_07249_),
    .Y(_07504_));
 sky130_fd_sc_hd__xnor2_1 _14334_ (.A(_07484_),
    .B(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__o22a_1 _14335_ (.A1(_07423_),
    .A2(_07303_),
    .B1(_07398_),
    .B2(_06959_),
    .X(_07506_));
 sky130_fd_sc_hd__or2_1 _14336_ (.A(_06982_),
    .B(_07366_),
    .X(_07507_));
 sky130_fd_sc_hd__or3_1 _14337_ (.A(_06757_),
    .B(_07417_),
    .C(_07366_),
    .X(_07508_));
 sky130_fd_sc_hd__a21oi_1 _14338_ (.A1(_07507_),
    .A2(_07508_),
    .B1(_07426_),
    .Y(_07509_));
 sky130_fd_sc_hd__a21oi_1 _14339_ (.A1(_07424_),
    .A2(_07506_),
    .B1(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__a21o_1 _14340_ (.A1(_07505_),
    .A2(_07510_),
    .B1(_07509_),
    .X(_07511_));
 sky130_fd_sc_hd__xnor2_1 _14341_ (.A(_07503_),
    .B(_07511_),
    .Y(_07512_));
 sky130_fd_sc_hd__and2b_1 _14342_ (.A_N(_07503_),
    .B(_07511_),
    .X(_07513_));
 sky130_fd_sc_hd__a21oi_1 _14343_ (.A1(_07500_),
    .A2(_07512_),
    .B1(_07513_),
    .Y(_07514_));
 sky130_fd_sc_hd__nor2_1 _14344_ (.A(_07499_),
    .B(_07514_),
    .Y(_07515_));
 sky130_fd_sc_hd__and2_1 _14345_ (.A(_07499_),
    .B(_07514_),
    .X(_07516_));
 sky130_fd_sc_hd__nor2_1 _14346_ (.A(_07515_),
    .B(_07516_),
    .Y(_07517_));
 sky130_fd_sc_hd__a21oi_1 _14347_ (.A1(_07498_),
    .A2(_07517_),
    .B1(_07515_),
    .Y(_07518_));
 sky130_fd_sc_hd__xnor2_1 _14348_ (.A(_07475_),
    .B(_07518_),
    .Y(_07519_));
 sky130_fd_sc_hd__nor2_1 _14349_ (.A(_07481_),
    .B(_07496_),
    .Y(_07520_));
 sky130_fd_sc_hd__a31o_1 _14350_ (.A1(_07446_),
    .A2(_07478_),
    .A3(_07497_),
    .B1(_07520_),
    .X(_07521_));
 sky130_fd_sc_hd__or2b_1 _14351_ (.A(_07519_),
    .B_N(_07521_),
    .X(_07522_));
 sky130_fd_sc_hd__o21a_1 _14352_ (.A1(_07475_),
    .A2(_07518_),
    .B1(_07522_),
    .X(_07523_));
 sky130_fd_sc_hd__nor2_1 _14353_ (.A(_07473_),
    .B(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__xor2_2 _14354_ (.A(_07413_),
    .B(_07466_),
    .X(_07525_));
 sky130_fd_sc_hd__and2_1 _14355_ (.A(_07524_),
    .B(_07525_),
    .X(_07526_));
 sky130_fd_sc_hd__and2_1 _14356_ (.A(_07472_),
    .B(_07526_),
    .X(_07527_));
 sky130_fd_sc_hd__nor2_1 _14357_ (.A(_07472_),
    .B(_07526_),
    .Y(_07528_));
 sky130_fd_sc_hd__nor2_1 _14358_ (.A(_07527_),
    .B(_07528_),
    .Y(_07529_));
 sky130_fd_sc_hd__inv_2 _14359_ (.A(_07529_),
    .Y(_07530_));
 sky130_fd_sc_hd__xor2_2 _14360_ (.A(_07521_),
    .B(_07519_),
    .X(_07531_));
 sky130_fd_sc_hd__or2_1 _14361_ (.A(_07045_),
    .B(_07248_),
    .X(_07532_));
 sky130_fd_sc_hd__or3b_1 _14362_ (.A(_07532_),
    .B(_07253_),
    .C_N(_07309_),
    .X(_07533_));
 sky130_fd_sc_hd__nor2_1 _14363_ (.A(_07253_),
    .B(_07248_),
    .Y(_07534_));
 sky130_fd_sc_hd__a21o_1 _14364_ (.A1(_06741_),
    .A2(_07310_),
    .B1(_07534_),
    .X(_07535_));
 sky130_fd_sc_hd__nor2_1 _14365_ (.A(_06942_),
    .B(_07204_),
    .Y(_07536_));
 sky130_fd_sc_hd__nand3_1 _14366_ (.A(_07533_),
    .B(_07535_),
    .C(_07536_),
    .Y(_07537_));
 sky130_fd_sc_hd__xnor2_1 _14367_ (.A(_07490_),
    .B(_07493_),
    .Y(_07538_));
 sky130_fd_sc_hd__a21oi_1 _14368_ (.A1(_07533_),
    .A2(_07537_),
    .B1(_07538_),
    .Y(_07539_));
 sky130_fd_sc_hd__and3_1 _14369_ (.A(_07533_),
    .B(_07537_),
    .C(_07538_),
    .X(_07540_));
 sky130_fd_sc_hd__or2_1 _14370_ (.A(_07539_),
    .B(_07540_),
    .X(_07541_));
 sky130_fd_sc_hd__or2_1 _14371_ (.A(_06993_),
    .B(_07360_),
    .X(_07542_));
 sky130_fd_sc_hd__inv_2 _14372_ (.A(_07542_),
    .Y(_07543_));
 sky130_fd_sc_hd__or2_1 _14373_ (.A(_07316_),
    .B(_07443_),
    .X(_07544_));
 sky130_fd_sc_hd__o21a_1 _14374_ (.A1(_07306_),
    .A2(_07361_),
    .B1(_07489_),
    .X(_07545_));
 sky130_fd_sc_hd__a21o_1 _14375_ (.A1(_07491_),
    .A2(_07543_),
    .B1(_07545_),
    .X(_07546_));
 sky130_fd_sc_hd__o2bb2a_1 _14376_ (.A1_N(_07491_),
    .A2_N(_07543_),
    .B1(_07544_),
    .B2(_07546_),
    .X(_07547_));
 sky130_fd_sc_hd__nor2_1 _14377_ (.A(_07541_),
    .B(_07547_),
    .Y(_07548_));
 sky130_fd_sc_hd__or2_1 _14378_ (.A(_07446_),
    .B(_07478_),
    .X(_07549_));
 sky130_fd_sc_hd__o211a_1 _14379_ (.A1(_07362_),
    .A2(_07445_),
    .B1(_07479_),
    .C1(_07549_),
    .X(_07550_));
 sky130_fd_sc_hd__o21a_1 _14380_ (.A1(_07539_),
    .A2(_07548_),
    .B1(_07550_),
    .X(_07551_));
 sky130_fd_sc_hd__xnor2_1 _14381_ (.A(_07498_),
    .B(_07517_),
    .Y(_07552_));
 sky130_fd_sc_hd__nor3_1 _14382_ (.A(_07539_),
    .B(_07548_),
    .C(_07550_),
    .Y(_07553_));
 sky130_fd_sc_hd__nor2_1 _14383_ (.A(_07551_),
    .B(_07553_),
    .Y(_07554_));
 sky130_fd_sc_hd__xnor2_1 _14384_ (.A(_07500_),
    .B(_07512_),
    .Y(_07555_));
 sky130_fd_sc_hd__xor2_1 _14385_ (.A(_07541_),
    .B(_07547_),
    .X(_07556_));
 sky130_fd_sc_hd__a21o_1 _14386_ (.A1(_07533_),
    .A2(_07535_),
    .B1(_07536_),
    .X(_07557_));
 sky130_fd_sc_hd__and2_1 _14387_ (.A(_07537_),
    .B(_07557_),
    .X(_07558_));
 sky130_fd_sc_hd__a21oi_1 _14388_ (.A1(_06757_),
    .A2(_07417_),
    .B1(_07303_),
    .Y(_07559_));
 sky130_fd_sc_hd__nand2_1 _14389_ (.A(_07508_),
    .B(_07559_),
    .Y(_07560_));
 sky130_fd_sc_hd__or4b_1 _14390_ (.A(_06757_),
    .B(_06785_),
    .C(_07366_),
    .D_N(_07309_),
    .X(_07561_));
 sky130_fd_sc_hd__nand2_1 _14391_ (.A(_07507_),
    .B(_07561_),
    .Y(_07562_));
 sky130_fd_sc_hd__xnor2_1 _14392_ (.A(_07560_),
    .B(_07562_),
    .Y(_07563_));
 sky130_fd_sc_hd__or2b_1 _14393_ (.A(_07560_),
    .B_N(_07562_),
    .X(_07564_));
 sky130_fd_sc_hd__a21bo_1 _14394_ (.A1(_07558_),
    .A2(_07563_),
    .B1_N(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__xnor2_1 _14395_ (.A(_07505_),
    .B(_07510_),
    .Y(_07566_));
 sky130_fd_sc_hd__xnor2_1 _14396_ (.A(_07565_),
    .B(_07566_),
    .Y(_07567_));
 sky130_fd_sc_hd__nand2_1 _14397_ (.A(_07558_),
    .B(_07563_),
    .Y(_07568_));
 sky130_fd_sc_hd__a21oi_1 _14398_ (.A1(_07564_),
    .A2(_07568_),
    .B1(_07566_),
    .Y(_07569_));
 sky130_fd_sc_hd__a21oi_1 _14399_ (.A1(_07556_),
    .A2(_07567_),
    .B1(_07569_),
    .Y(_07570_));
 sky130_fd_sc_hd__xor2_1 _14400_ (.A(_07555_),
    .B(_07570_),
    .X(_07571_));
 sky130_fd_sc_hd__nor2_1 _14401_ (.A(_07555_),
    .B(_07570_),
    .Y(_07572_));
 sky130_fd_sc_hd__a21oi_1 _14402_ (.A1(_07554_),
    .A2(_07571_),
    .B1(_07572_),
    .Y(_07573_));
 sky130_fd_sc_hd__xor2_1 _14403_ (.A(_07552_),
    .B(_07573_),
    .X(_07574_));
 sky130_fd_sc_hd__nor2_1 _14404_ (.A(_07552_),
    .B(_07573_),
    .Y(_07575_));
 sky130_fd_sc_hd__a21oi_2 _14405_ (.A1(_07551_),
    .A2(_07574_),
    .B1(_07575_),
    .Y(_07576_));
 sky130_fd_sc_hd__nor2_1 _14406_ (.A(_07531_),
    .B(_07576_),
    .Y(_07577_));
 sky130_fd_sc_hd__xor2_2 _14407_ (.A(_07473_),
    .B(_07523_),
    .X(_07578_));
 sky130_fd_sc_hd__and2_1 _14408_ (.A(_07577_),
    .B(_07578_),
    .X(_07579_));
 sky130_fd_sc_hd__xnor2_1 _14409_ (.A(_07551_),
    .B(_07574_),
    .Y(_07580_));
 sky130_fd_sc_hd__nor2_1 _14410_ (.A(_07045_),
    .B(_07204_),
    .Y(_07581_));
 sky130_fd_sc_hd__nand2_1 _14411_ (.A(_07534_),
    .B(_07581_),
    .Y(_07582_));
 sky130_fd_sc_hd__nor2_1 _14412_ (.A(_07253_),
    .B(_07204_),
    .Y(_07583_));
 sky130_fd_sc_hd__xnor2_1 _14413_ (.A(_07532_),
    .B(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__nor2_1 _14414_ (.A(_06942_),
    .B(_07209_),
    .Y(_07585_));
 sky130_fd_sc_hd__nand2_1 _14415_ (.A(_07584_),
    .B(_07585_),
    .Y(_07586_));
 sky130_fd_sc_hd__xnor2_1 _14416_ (.A(_07544_),
    .B(_07546_),
    .Y(_07587_));
 sky130_fd_sc_hd__a21o_1 _14417_ (.A1(_07582_),
    .A2(_07586_),
    .B1(_07587_),
    .X(_07588_));
 sky130_fd_sc_hd__nand3_1 _14418_ (.A(_07582_),
    .B(_07586_),
    .C(_07587_),
    .Y(_07589_));
 sky130_fd_sc_hd__nand2_1 _14419_ (.A(_07588_),
    .B(_07589_),
    .Y(_07590_));
 sky130_fd_sc_hd__nor2_1 _14420_ (.A(_07306_),
    .B(_07443_),
    .Y(_07591_));
 sky130_fd_sc_hd__inv_2 _14421_ (.A(_07591_),
    .Y(_07592_));
 sky130_fd_sc_hd__xnor2_1 _14422_ (.A(_07542_),
    .B(_07592_),
    .Y(_07593_));
 sky130_fd_sc_hd__o32a_1 _14423_ (.A1(_07316_),
    .A2(_07476_),
    .A3(_07593_),
    .B1(_07592_),
    .B2(_07542_),
    .X(_07594_));
 sky130_fd_sc_hd__or2_1 _14424_ (.A(_07590_),
    .B(_07594_),
    .X(_07595_));
 sky130_fd_sc_hd__o22a_1 _14425_ (.A1(_07206_),
    .A2(_07476_),
    .B1(_07444_),
    .B2(_06720_),
    .X(_07596_));
 sky130_fd_sc_hd__or2_1 _14426_ (.A(_07478_),
    .B(_07596_),
    .X(_07597_));
 sky130_fd_sc_hd__a21oi_2 _14427_ (.A1(_07588_),
    .A2(_07595_),
    .B1(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__xnor2_1 _14428_ (.A(_07554_),
    .B(_07571_),
    .Y(_07599_));
 sky130_fd_sc_hd__and3_1 _14429_ (.A(_07588_),
    .B(_07595_),
    .C(_07597_),
    .X(_07600_));
 sky130_fd_sc_hd__nor2_1 _14430_ (.A(_07598_),
    .B(_07600_),
    .Y(_07601_));
 sky130_fd_sc_hd__xnor2_1 _14431_ (.A(_07556_),
    .B(_07567_),
    .Y(_07602_));
 sky130_fd_sc_hd__xor2_1 _14432_ (.A(_07590_),
    .B(_07594_),
    .X(_07603_));
 sky130_fd_sc_hd__xnor2_1 _14433_ (.A(_07558_),
    .B(_07563_),
    .Y(_07604_));
 sky130_fd_sc_hd__or2_1 _14434_ (.A(_07584_),
    .B(_07585_),
    .X(_07605_));
 sky130_fd_sc_hd__and2_1 _14435_ (.A(_07586_),
    .B(_07605_),
    .X(_07606_));
 sky130_fd_sc_hd__a2bb2o_1 _14436_ (.A1_N(_06757_),
    .A2_N(_07303_),
    .B1(_07310_),
    .B2(_06807_),
    .X(_07607_));
 sky130_fd_sc_hd__nand2_1 _14437_ (.A(_07561_),
    .B(_07607_),
    .Y(_07608_));
 sky130_fd_sc_hd__nor2_1 _14438_ (.A(_07417_),
    .B(_07248_),
    .Y(_07609_));
 sky130_fd_sc_hd__a2bb2o_1 _14439_ (.A1_N(_06959_),
    .A2_N(_07366_),
    .B1(_07310_),
    .B2(_06808_),
    .X(_07610_));
 sky130_fd_sc_hd__or4b_1 _14440_ (.A(_06959_),
    .B(_07423_),
    .C(_07366_),
    .D_N(_07309_),
    .X(_07611_));
 sky130_fd_sc_hd__a21boi_1 _14441_ (.A1(_07609_),
    .A2(_07610_),
    .B1_N(_07611_),
    .Y(_07612_));
 sky130_fd_sc_hd__xor2_1 _14442_ (.A(_07608_),
    .B(_07612_),
    .X(_07613_));
 sky130_fd_sc_hd__nor2_1 _14443_ (.A(_07608_),
    .B(_07612_),
    .Y(_07614_));
 sky130_fd_sc_hd__a21oi_1 _14444_ (.A1(_07606_),
    .A2(_07613_),
    .B1(_07614_),
    .Y(_07615_));
 sky130_fd_sc_hd__xor2_1 _14445_ (.A(_07604_),
    .B(_07615_),
    .X(_07616_));
 sky130_fd_sc_hd__nor2_1 _14446_ (.A(_07604_),
    .B(_07615_),
    .Y(_07617_));
 sky130_fd_sc_hd__a21oi_1 _14447_ (.A1(_07603_),
    .A2(_07616_),
    .B1(_07617_),
    .Y(_07618_));
 sky130_fd_sc_hd__xor2_1 _14448_ (.A(_07602_),
    .B(_07618_),
    .X(_07619_));
 sky130_fd_sc_hd__nor2_1 _14449_ (.A(_07602_),
    .B(_07618_),
    .Y(_07620_));
 sky130_fd_sc_hd__a21oi_1 _14450_ (.A1(_07601_),
    .A2(_07619_),
    .B1(_07620_),
    .Y(_07621_));
 sky130_fd_sc_hd__xor2_1 _14451_ (.A(_07599_),
    .B(_07621_),
    .X(_07622_));
 sky130_fd_sc_hd__nor2_1 _14452_ (.A(_07599_),
    .B(_07621_),
    .Y(_07623_));
 sky130_fd_sc_hd__a21oi_2 _14453_ (.A1(_07598_),
    .A2(_07622_),
    .B1(_07623_),
    .Y(_07624_));
 sky130_fd_sc_hd__nor2_1 _14454_ (.A(_07580_),
    .B(_07624_),
    .Y(_07625_));
 sky130_fd_sc_hd__xor2_2 _14455_ (.A(_07531_),
    .B(_07576_),
    .X(_07626_));
 sky130_fd_sc_hd__and2_1 _14456_ (.A(_07625_),
    .B(_07626_),
    .X(_07627_));
 sky130_fd_sc_hd__xnor2_1 _14457_ (.A(_07598_),
    .B(_07622_),
    .Y(_07628_));
 sky130_fd_sc_hd__nor2_1 _14458_ (.A(_06857_),
    .B(_07209_),
    .Y(_07629_));
 sky130_fd_sc_hd__nand2_1 _14459_ (.A(_07581_),
    .B(_07629_),
    .Y(_07630_));
 sky130_fd_sc_hd__or2_1 _14460_ (.A(_07581_),
    .B(_07629_),
    .X(_07631_));
 sky130_fd_sc_hd__nand2_1 _14461_ (.A(_07630_),
    .B(_07631_),
    .Y(_07632_));
 sky130_fd_sc_hd__or3_1 _14462_ (.A(_07252_),
    .B(_07361_),
    .C(_07632_),
    .X(_07633_));
 sky130_fd_sc_hd__or2_1 _14463_ (.A(_07316_),
    .B(_07158_),
    .X(_07634_));
 sky130_fd_sc_hd__xnor2_1 _14464_ (.A(_07634_),
    .B(_07593_),
    .Y(_07635_));
 sky130_fd_sc_hd__a21o_1 _14465_ (.A1(_07630_),
    .A2(_07633_),
    .B1(_07635_),
    .X(_07636_));
 sky130_fd_sc_hd__nand3_1 _14466_ (.A(_07630_),
    .B(_07633_),
    .C(_07635_),
    .Y(_07637_));
 sky130_fd_sc_hd__nand2_1 _14467_ (.A(_07636_),
    .B(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__or2_1 _14468_ (.A(_06993_),
    .B(_07476_),
    .X(_07639_));
 sky130_fd_sc_hd__clkbuf_2 _14469_ (.A(_07639_),
    .X(_07640_));
 sky130_fd_sc_hd__o31a_1 _14470_ (.A1(_07592_),
    .A2(_07638_),
    .A3(_07640_),
    .B1(_07636_),
    .X(_07641_));
 sky130_fd_sc_hd__nor2b_1 _14471_ (.A(_07641_),
    .B_N(_07477_),
    .Y(_07642_));
 sky130_fd_sc_hd__xnor2_1 _14472_ (.A(_07601_),
    .B(_07619_),
    .Y(_07643_));
 sky130_fd_sc_hd__and2b_1 _14473_ (.A_N(_07477_),
    .B(_07641_),
    .X(_07644_));
 sky130_fd_sc_hd__nor2_1 _14474_ (.A(_07642_),
    .B(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__xnor2_1 _14475_ (.A(_07603_),
    .B(_07616_),
    .Y(_07646_));
 sky130_fd_sc_hd__nor2_1 _14476_ (.A(_07592_),
    .B(_07640_),
    .Y(_07647_));
 sky130_fd_sc_hd__xnor2_1 _14477_ (.A(_07638_),
    .B(_07647_),
    .Y(_07648_));
 sky130_fd_sc_hd__xnor2_1 _14478_ (.A(_07606_),
    .B(_07613_),
    .Y(_07649_));
 sky130_fd_sc_hd__nor2_1 _14479_ (.A(_07252_),
    .B(_07361_),
    .Y(_07650_));
 sky130_fd_sc_hd__xnor2_1 _14480_ (.A(_07632_),
    .B(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__nand3_1 _14481_ (.A(_07611_),
    .B(_07609_),
    .C(_07610_),
    .Y(_07652_));
 sky130_fd_sc_hd__a21o_1 _14482_ (.A1(_07611_),
    .A2(_07610_),
    .B1(_07609_),
    .X(_07653_));
 sky130_fd_sc_hd__nor2_1 _14483_ (.A(_07417_),
    .B(_07204_),
    .Y(_07654_));
 sky130_fd_sc_hd__nor2_1 _14484_ (.A(_07423_),
    .B(_07248_),
    .Y(_07655_));
 sky130_fd_sc_hd__a21o_1 _14485_ (.A1(_06729_),
    .A2(_07310_),
    .B1(_07655_),
    .X(_07656_));
 sky130_fd_sc_hd__nand3_1 _14486_ (.A(_06729_),
    .B(_07310_),
    .C(_07655_),
    .Y(_07657_));
 sky130_fd_sc_hd__a21bo_1 _14487_ (.A1(_07654_),
    .A2(_07656_),
    .B1_N(_07657_),
    .X(_07658_));
 sky130_fd_sc_hd__a21o_1 _14488_ (.A1(_07652_),
    .A2(_07653_),
    .B1(_07658_),
    .X(_07659_));
 sky130_fd_sc_hd__nand3_1 _14489_ (.A(_07652_),
    .B(_07653_),
    .C(_07658_),
    .Y(_07660_));
 sky130_fd_sc_hd__a21boi_1 _14490_ (.A1(_07651_),
    .A2(_07659_),
    .B1_N(_07660_),
    .Y(_07661_));
 sky130_fd_sc_hd__xor2_1 _14491_ (.A(_07649_),
    .B(_07661_),
    .X(_07662_));
 sky130_fd_sc_hd__nor2_1 _14492_ (.A(_07649_),
    .B(_07661_),
    .Y(_07663_));
 sky130_fd_sc_hd__a21o_1 _14493_ (.A1(_07648_),
    .A2(_07662_),
    .B1(_07663_),
    .X(_07664_));
 sky130_fd_sc_hd__xnor2_1 _14494_ (.A(_07646_),
    .B(_07664_),
    .Y(_07665_));
 sky130_fd_sc_hd__or2b_1 _14495_ (.A(_07646_),
    .B_N(_07664_),
    .X(_07666_));
 sky130_fd_sc_hd__a21boi_1 _14496_ (.A1(_07645_),
    .A2(_07665_),
    .B1_N(_07666_),
    .Y(_07667_));
 sky130_fd_sc_hd__xor2_1 _14497_ (.A(_07643_),
    .B(_07667_),
    .X(_07668_));
 sky130_fd_sc_hd__nor2_1 _14498_ (.A(_07643_),
    .B(_07667_),
    .Y(_07669_));
 sky130_fd_sc_hd__a21oi_2 _14499_ (.A1(_07642_),
    .A2(_07668_),
    .B1(_07669_),
    .Y(_07670_));
 sky130_fd_sc_hd__nor2_1 _14500_ (.A(_07628_),
    .B(_07670_),
    .Y(_07671_));
 sky130_fd_sc_hd__xor2_1 _14501_ (.A(_07580_),
    .B(_07624_),
    .X(_07672_));
 sky130_fd_sc_hd__and2_1 _14502_ (.A(_07671_),
    .B(_07672_),
    .X(_07673_));
 sky130_fd_sc_hd__xor2_1 _14503_ (.A(_07628_),
    .B(_07670_),
    .X(_07674_));
 sky130_fd_sc_hd__nor2_1 _14504_ (.A(_07045_),
    .B(_07361_),
    .Y(_07675_));
 sky130_fd_sc_hd__nand2_1 _14505_ (.A(_07629_),
    .B(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__o22a_1 _14506_ (.A1(_07045_),
    .A2(_07209_),
    .B1(_07361_),
    .B2(_07253_),
    .X(_07677_));
 sky130_fd_sc_hd__a21o_1 _14507_ (.A1(_07629_),
    .A2(_07675_),
    .B1(_07677_),
    .X(_07678_));
 sky130_fd_sc_hd__or3_1 _14508_ (.A(_07252_),
    .B(_07444_),
    .C(_07678_),
    .X(_07679_));
 sky130_fd_sc_hd__o22a_1 _14509_ (.A1(_07306_),
    .A2(_07476_),
    .B1(_07444_),
    .B2(_06993_),
    .X(_07680_));
 sky130_fd_sc_hd__or2_1 _14510_ (.A(_07647_),
    .B(_07680_),
    .X(_07681_));
 sky130_fd_sc_hd__a21oi_2 _14511_ (.A1(_07676_),
    .A2(_07679_),
    .B1(_07681_),
    .Y(_07682_));
 sky130_fd_sc_hd__xnor2_1 _14512_ (.A(_07648_),
    .B(_07662_),
    .Y(_07683_));
 sky130_fd_sc_hd__and3_1 _14513_ (.A(_07676_),
    .B(_07679_),
    .C(_07681_),
    .X(_07684_));
 sky130_fd_sc_hd__nor2_1 _14514_ (.A(_07682_),
    .B(_07684_),
    .Y(_07685_));
 sky130_fd_sc_hd__nand3_1 _14515_ (.A(_07660_),
    .B(_07651_),
    .C(_07659_),
    .Y(_07686_));
 sky130_fd_sc_hd__a21o_1 _14516_ (.A1(_07660_),
    .A2(_07659_),
    .B1(_07651_),
    .X(_07687_));
 sky130_fd_sc_hd__nor2_1 _14517_ (.A(_07252_),
    .B(_07444_),
    .Y(_07688_));
 sky130_fd_sc_hd__xnor2_1 _14518_ (.A(_07678_),
    .B(_07688_),
    .Y(_07689_));
 sky130_fd_sc_hd__nand3_1 _14519_ (.A(_07657_),
    .B(_07654_),
    .C(_07656_),
    .Y(_07690_));
 sky130_fd_sc_hd__a21o_1 _14520_ (.A1(_07657_),
    .A2(_07656_),
    .B1(_07654_),
    .X(_07691_));
 sky130_fd_sc_hd__or2_1 _14521_ (.A(_06959_),
    .B(_07204_),
    .X(_07692_));
 sky130_fd_sc_hd__nor3_1 _14522_ (.A(_07423_),
    .B(_07248_),
    .C(_07692_),
    .Y(_07693_));
 sky130_fd_sc_hd__nor2_1 _14523_ (.A(_07417_),
    .B(_07209_),
    .Y(_07694_));
 sky130_fd_sc_hd__inv_2 _14524_ (.A(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__nor2_1 _14525_ (.A(_07423_),
    .B(_07204_),
    .Y(_07696_));
 sky130_fd_sc_hd__o21ba_1 _14526_ (.A1(_06959_),
    .A2(_07248_),
    .B1_N(_07696_),
    .X(_07697_));
 sky130_fd_sc_hd__or3_2 _14527_ (.A(_07693_),
    .B(_07695_),
    .C(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__or2b_1 _14528_ (.A(_07693_),
    .B_N(_07698_),
    .X(_07699_));
 sky130_fd_sc_hd__a21o_1 _14529_ (.A1(_07690_),
    .A2(_07691_),
    .B1(_07699_),
    .X(_07700_));
 sky130_fd_sc_hd__nand3_1 _14530_ (.A(_07690_),
    .B(_07691_),
    .C(_07699_),
    .Y(_07701_));
 sky130_fd_sc_hd__a21bo_1 _14531_ (.A1(_07689_),
    .A2(_07700_),
    .B1_N(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__and3_1 _14532_ (.A(_07686_),
    .B(_07687_),
    .C(_07702_),
    .X(_07703_));
 sky130_fd_sc_hd__a21oi_1 _14533_ (.A1(_07686_),
    .A2(_07687_),
    .B1(_07702_),
    .Y(_07704_));
 sky130_fd_sc_hd__nor2_1 _14534_ (.A(_07703_),
    .B(_07704_),
    .Y(_07705_));
 sky130_fd_sc_hd__a21oi_1 _14535_ (.A1(_07685_),
    .A2(_07705_),
    .B1(_07703_),
    .Y(_07706_));
 sky130_fd_sc_hd__nand2_1 _14536_ (.A(_07683_),
    .B(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__nor2_1 _14537_ (.A(_07683_),
    .B(_07706_),
    .Y(_07708_));
 sky130_fd_sc_hd__a21oi_2 _14538_ (.A1(_07682_),
    .A2(_07707_),
    .B1(_07708_),
    .Y(_07709_));
 sky130_fd_sc_hd__xnor2_1 _14539_ (.A(_07645_),
    .B(_07665_),
    .Y(_07710_));
 sky130_fd_sc_hd__xor2_1 _14540_ (.A(_07642_),
    .B(_07668_),
    .X(_07711_));
 sky130_fd_sc_hd__nor3b_2 _14541_ (.A(_07709_),
    .B(_07710_),
    .C_N(_07711_),
    .Y(_07712_));
 sky130_fd_sc_hd__and2_1 _14542_ (.A(_07674_),
    .B(_07712_),
    .X(_07713_));
 sky130_fd_sc_hd__xor2_1 _14543_ (.A(_07674_),
    .B(_07712_),
    .X(_07714_));
 sky130_fd_sc_hd__and2b_1 _14544_ (.A_N(_07708_),
    .B(_07707_),
    .X(_07715_));
 sky130_fd_sc_hd__xor2_1 _14545_ (.A(_07682_),
    .B(_07715_),
    .X(_07716_));
 sky130_fd_sc_hd__xnor2_1 _14546_ (.A(_07685_),
    .B(_07705_),
    .Y(_07717_));
 sky130_fd_sc_hd__nor2_1 _14547_ (.A(_07253_),
    .B(_07444_),
    .Y(_07718_));
 sky130_fd_sc_hd__nand2_1 _14548_ (.A(_07675_),
    .B(_07718_),
    .Y(_07719_));
 sky130_fd_sc_hd__or2_1 _14549_ (.A(_07675_),
    .B(_07718_),
    .X(_07720_));
 sky130_fd_sc_hd__nand2_1 _14550_ (.A(_07719_),
    .B(_07720_),
    .Y(_07721_));
 sky130_fd_sc_hd__o31a_1 _14551_ (.A1(_07252_),
    .A2(_07476_),
    .A3(_07721_),
    .B1(_07719_),
    .X(_07722_));
 sky130_fd_sc_hd__xor2_1 _14552_ (.A(_07640_),
    .B(_07722_),
    .X(_07723_));
 sky130_fd_sc_hd__nand2_1 _14553_ (.A(_07701_),
    .B(_07700_),
    .Y(_07724_));
 sky130_fd_sc_hd__xor2_1 _14554_ (.A(_07689_),
    .B(_07724_),
    .X(_07725_));
 sky130_fd_sc_hd__o21ai_2 _14555_ (.A1(_07693_),
    .A2(_07697_),
    .B1(_07695_),
    .Y(_07726_));
 sky130_fd_sc_hd__nor2_1 _14556_ (.A(_06959_),
    .B(_07209_),
    .Y(_07727_));
 sky130_fd_sc_hd__nor2_1 _14557_ (.A(_07417_),
    .B(_07361_),
    .Y(_07728_));
 sky130_fd_sc_hd__nor2_1 _14558_ (.A(_07423_),
    .B(_07209_),
    .Y(_07729_));
 sky130_fd_sc_hd__xnor2_1 _14559_ (.A(_07692_),
    .B(_07729_),
    .Y(_07730_));
 sky130_fd_sc_hd__a22o_2 _14560_ (.A1(_07696_),
    .A2(_07727_),
    .B1(_07728_),
    .B2(_07730_),
    .X(_07731_));
 sky130_fd_sc_hd__nor2_1 _14561_ (.A(_07252_),
    .B(_07476_),
    .Y(_07732_));
 sky130_fd_sc_hd__xnor2_2 _14562_ (.A(_07721_),
    .B(_07732_),
    .Y(_07733_));
 sky130_fd_sc_hd__nand2_1 _14563_ (.A(_07698_),
    .B(_07726_),
    .Y(_07734_));
 sky130_fd_sc_hd__xnor2_2 _14564_ (.A(_07734_),
    .B(_07731_),
    .Y(_07735_));
 sky130_fd_sc_hd__a32oi_4 _14565_ (.A1(_07698_),
    .A2(_07726_),
    .A3(_07731_),
    .B1(_07733_),
    .B2(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__xor2_1 _14566_ (.A(_07725_),
    .B(_07736_),
    .X(_07737_));
 sky130_fd_sc_hd__nor2_1 _14567_ (.A(_07725_),
    .B(_07736_),
    .Y(_07738_));
 sky130_fd_sc_hd__a21oi_1 _14568_ (.A1(_07723_),
    .A2(_07737_),
    .B1(_07738_),
    .Y(_07739_));
 sky130_fd_sc_hd__xnor2_1 _14569_ (.A(_07717_),
    .B(_07739_),
    .Y(_07740_));
 sky130_fd_sc_hd__nor3_1 _14570_ (.A(_07640_),
    .B(_07722_),
    .C(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__o21bai_1 _14571_ (.A1(_07717_),
    .A2(_07739_),
    .B1_N(_07741_),
    .Y(_07742_));
 sky130_fd_sc_hd__xor2_1 _14572_ (.A(_07710_),
    .B(_07709_),
    .X(_07743_));
 sky130_fd_sc_hd__and4_1 _14573_ (.A(_07711_),
    .B(_07716_),
    .C(_07742_),
    .D(_07743_),
    .X(_07744_));
 sky130_fd_sc_hd__xor2_1 _14574_ (.A(_07714_),
    .B(_07744_),
    .X(_07745_));
 sky130_fd_sc_hd__nand2_1 _14575_ (.A(_07711_),
    .B(_07743_),
    .Y(_07746_));
 sky130_fd_sc_hd__nor2_1 _14576_ (.A(_07716_),
    .B(_07742_),
    .Y(_07747_));
 sky130_fd_sc_hd__o21a_1 _14577_ (.A1(_07640_),
    .A2(_07722_),
    .B1(_07740_),
    .X(_07748_));
 sky130_fd_sc_hd__nor2_1 _14578_ (.A(_07417_),
    .B(_07444_),
    .Y(_07749_));
 sky130_fd_sc_hd__nor2_1 _14579_ (.A(_07423_),
    .B(_07361_),
    .Y(_07750_));
 sky130_fd_sc_hd__xor2_1 _14580_ (.A(_07727_),
    .B(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__xor2_1 _14581_ (.A(_07749_),
    .B(_07751_),
    .X(_07752_));
 sky130_fd_sc_hd__inv_2 _14582_ (.A(_07752_),
    .Y(_07753_));
 sky130_fd_sc_hd__or2_1 _14583_ (.A(_06959_),
    .B(_07361_),
    .X(_07754_));
 sky130_fd_sc_hd__nor2_1 _14584_ (.A(_07417_),
    .B(_07476_),
    .Y(_07755_));
 sky130_fd_sc_hd__nor2_1 _14585_ (.A(_07423_),
    .B(_07444_),
    .Y(_07756_));
 sky130_fd_sc_hd__xnor2_1 _14586_ (.A(_07754_),
    .B(_07756_),
    .Y(_07757_));
 sky130_fd_sc_hd__nand2_1 _14587_ (.A(_07755_),
    .B(_07757_),
    .Y(_07758_));
 sky130_fd_sc_hd__o31a_1 _14588_ (.A1(_07423_),
    .A2(_07444_),
    .A3(_07754_),
    .B1(_07758_),
    .X(_07759_));
 sky130_fd_sc_hd__nor2_1 _14589_ (.A(_07045_),
    .B(_07476_),
    .Y(_07760_));
 sky130_fd_sc_hd__xnor2_1 _14590_ (.A(_07752_),
    .B(_07759_),
    .Y(_07761_));
 sky130_fd_sc_hd__nand2_1 _14591_ (.A(_07760_),
    .B(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__o21ai_1 _14592_ (.A1(_07753_),
    .A2(_07759_),
    .B1(_07762_),
    .Y(_07763_));
 sky130_fd_sc_hd__or2_1 _14593_ (.A(_07760_),
    .B(_07761_),
    .X(_07764_));
 sky130_fd_sc_hd__and3b_1 _14594_ (.A_N(_06982_),
    .B(_07159_),
    .C(_07758_),
    .X(_07765_));
 sky130_fd_sc_hd__o2111a_1 _14595_ (.A1(_07755_),
    .A2(_07757_),
    .B1(_07762_),
    .C1(_07764_),
    .D1(_07765_),
    .X(_07766_));
 sky130_fd_sc_hd__nand2_1 _14596_ (.A(_07763_),
    .B(_07766_),
    .Y(_07767_));
 sky130_fd_sc_hd__and2_1 _14597_ (.A(_07718_),
    .B(_07760_),
    .X(_07768_));
 sky130_fd_sc_hd__o22a_1 _14598_ (.A1(_07253_),
    .A2(_07476_),
    .B1(_07444_),
    .B2(_07045_),
    .X(_07769_));
 sky130_fd_sc_hd__nor2_1 _14599_ (.A(_07768_),
    .B(_07769_),
    .Y(_07770_));
 sky130_fd_sc_hd__xnor2_1 _14600_ (.A(_07728_),
    .B(_07730_),
    .Y(_07771_));
 sky130_fd_sc_hd__a22oi_1 _14601_ (.A1(_07727_),
    .A2(_07750_),
    .B1(_07749_),
    .B2(_07751_),
    .Y(_07772_));
 sky130_fd_sc_hd__or2_1 _14602_ (.A(_07771_),
    .B(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__nand2_1 _14603_ (.A(_07771_),
    .B(_07772_),
    .Y(_07774_));
 sky130_fd_sc_hd__and2_1 _14604_ (.A(_07773_),
    .B(_07774_),
    .X(_07775_));
 sky130_fd_sc_hd__nand2_1 _14605_ (.A(_07770_),
    .B(_07775_),
    .Y(_07776_));
 sky130_fd_sc_hd__or2_1 _14606_ (.A(_07770_),
    .B(_07775_),
    .X(_07777_));
 sky130_fd_sc_hd__nand2_1 _14607_ (.A(_07776_),
    .B(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__nor2_1 _14608_ (.A(_07763_),
    .B(_07766_),
    .Y(_07779_));
 sky130_fd_sc_hd__a21oi_1 _14609_ (.A1(_07767_),
    .A2(_07778_),
    .B1(_07779_),
    .Y(_07780_));
 sky130_fd_sc_hd__xnor2_1 _14610_ (.A(_07733_),
    .B(_07735_),
    .Y(_07781_));
 sky130_fd_sc_hd__and2_1 _14611_ (.A(_07773_),
    .B(_07776_),
    .X(_07782_));
 sky130_fd_sc_hd__a2bb2o_1 _14612_ (.A1_N(_07780_),
    .A2_N(_07768_),
    .B1(_07781_),
    .B2(_07782_),
    .X(_07783_));
 sky130_fd_sc_hd__o2bb2a_1 _14613_ (.A1_N(_07780_),
    .A2_N(_07768_),
    .B1(_07781_),
    .B2(_07782_),
    .X(_07784_));
 sky130_fd_sc_hd__nor2_1 _14614_ (.A(_07723_),
    .B(_07737_),
    .Y(_07785_));
 sky130_fd_sc_hd__a221oi_1 _14615_ (.A1(_07723_),
    .A2(_07737_),
    .B1(_07783_),
    .B2(_07784_),
    .C1(_07785_),
    .Y(_07786_));
 sky130_fd_sc_hd__or4b_1 _14616_ (.A(_07741_),
    .B(_07747_),
    .C(_07748_),
    .D_N(_07786_),
    .X(_07787_));
 sky130_fd_sc_hd__nor2_2 _14617_ (.A(_07746_),
    .B(_07787_),
    .Y(_07788_));
 sky130_fd_sc_hd__and2_1 _14618_ (.A(_07714_),
    .B(_07744_),
    .X(_07789_));
 sky130_fd_sc_hd__a21o_1 _14619_ (.A1(_07745_),
    .A2(_07788_),
    .B1(_07789_),
    .X(_07790_));
 sky130_fd_sc_hd__nor2_1 _14620_ (.A(_07671_),
    .B(_07713_),
    .Y(_07791_));
 sky130_fd_sc_hd__xnor2_1 _14621_ (.A(_07672_),
    .B(_07791_),
    .Y(_07792_));
 sky130_fd_sc_hd__a22o_1 _14622_ (.A1(_07713_),
    .A2(_07672_),
    .B1(_07790_),
    .B2(_07792_),
    .X(_07793_));
 sky130_fd_sc_hd__nor2_1 _14623_ (.A(_07625_),
    .B(_07673_),
    .Y(_07794_));
 sky130_fd_sc_hd__xnor2_1 _14624_ (.A(_07626_),
    .B(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__a22o_1 _14625_ (.A1(_07626_),
    .A2(_07673_),
    .B1(_07793_),
    .B2(_07795_),
    .X(_07796_));
 sky130_fd_sc_hd__nor3_1 _14626_ (.A(_07577_),
    .B(_07578_),
    .C(_07627_),
    .Y(_07797_));
 sky130_fd_sc_hd__a211oi_1 _14627_ (.A1(_07578_),
    .A2(_07627_),
    .B1(_07797_),
    .C1(_07579_),
    .Y(_07798_));
 sky130_fd_sc_hd__a22o_1 _14628_ (.A1(_07578_),
    .A2(_07627_),
    .B1(_07796_),
    .B2(_07798_),
    .X(_07799_));
 sky130_fd_sc_hd__nor2_1 _14629_ (.A(_07524_),
    .B(_07579_),
    .Y(_07800_));
 sky130_fd_sc_hd__xnor2_1 _14630_ (.A(_07525_),
    .B(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__a22oi_2 _14631_ (.A1(_07525_),
    .A2(_07579_),
    .B1(_07799_),
    .B2(_07801_),
    .Y(_07802_));
 sky130_fd_sc_hd__o21ba_1 _14632_ (.A1(_07530_),
    .A2(_07802_),
    .B1_N(_07527_),
    .X(_07803_));
 sky130_fd_sc_hd__xnor2_1 _14633_ (.A(_07471_),
    .B(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__xnor2_1 _14634_ (.A(_07529_),
    .B(_07802_),
    .Y(_07805_));
 sky130_fd_sc_hd__buf_2 _14635_ (.A(_06579_),
    .X(_07806_));
 sky130_fd_sc_hd__mux2_1 _14636_ (.A0(_07804_),
    .A1(_07805_),
    .S(_07806_),
    .X(_07807_));
 sky130_fd_sc_hd__xnor2_1 _14637_ (.A(_07796_),
    .B(_07798_),
    .Y(_07808_));
 sky130_fd_sc_hd__xnor2_1 _14638_ (.A(_07799_),
    .B(_07801_),
    .Y(_07809_));
 sky130_fd_sc_hd__nor2_1 _14639_ (.A(_06579_),
    .B(_07809_),
    .Y(_07810_));
 sky130_fd_sc_hd__o21ba_1 _14640_ (.A1(_06613_),
    .A2(_07808_),
    .B1_N(_07810_),
    .X(_07811_));
 sky130_fd_sc_hd__nand2_1 _14641_ (.A(_06580_),
    .B(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__o21ai_1 _14642_ (.A1(_06580_),
    .A2(_07807_),
    .B1(_07812_),
    .Y(_07813_));
 sky130_fd_sc_hd__xnor2_1 _14643_ (.A(_07745_),
    .B(_07788_),
    .Y(_07814_));
 sky130_fd_sc_hd__or2_1 _14644_ (.A(_07806_),
    .B(_07814_),
    .X(_07815_));
 sky130_fd_sc_hd__clkinv_2 _14645_ (.A(_07815_),
    .Y(_07816_));
 sky130_fd_sc_hd__xnor2_1 _14646_ (.A(_07793_),
    .B(_07795_),
    .Y(_07817_));
 sky130_fd_sc_hd__or2_1 _14647_ (.A(_06579_),
    .B(_07817_),
    .X(_07818_));
 sky130_fd_sc_hd__xnor2_1 _14648_ (.A(_07790_),
    .B(_07792_),
    .Y(_07819_));
 sky130_fd_sc_hd__or2_1 _14649_ (.A(_06613_),
    .B(_07819_),
    .X(_07820_));
 sky130_fd_sc_hd__nand2_1 _14650_ (.A(_07818_),
    .B(_07820_),
    .Y(_07821_));
 sky130_fd_sc_hd__buf_2 _14651_ (.A(_06584_),
    .X(_07822_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(_07816_),
    .A1(_07821_),
    .S(_07822_),
    .X(_07823_));
 sky130_fd_sc_hd__nand2_1 _14653_ (.A(_06574_),
    .B(_07823_),
    .Y(_07824_));
 sky130_fd_sc_hd__o21a_1 _14654_ (.A1(_06575_),
    .A2(_07813_),
    .B1(_07824_),
    .X(_07825_));
 sky130_fd_sc_hd__buf_2 _14655_ (.A(_06595_),
    .X(_07826_));
 sky130_fd_sc_hd__buf_2 _14656_ (.A(_06613_),
    .X(_07827_));
 sky130_fd_sc_hd__and2_1 _14657_ (.A(_06758_),
    .B(_07331_),
    .X(_07828_));
 sky130_fd_sc_hd__a21oi_1 _14658_ (.A1(_06758_),
    .A2(_06738_),
    .B1(_07331_),
    .Y(_07829_));
 sky130_fd_sc_hd__and2_1 _14659_ (.A(_07333_),
    .B(_07401_),
    .X(_07830_));
 sky130_fd_sc_hd__o21a_1 _14660_ (.A1(_07828_),
    .A2(_07829_),
    .B1(_07830_),
    .X(_07831_));
 sky130_fd_sc_hd__xnor2_1 _14661_ (.A(_07402_),
    .B(_07831_),
    .Y(_07832_));
 sky130_fd_sc_hd__xnor2_1 _14662_ (.A(_07407_),
    .B(_07832_),
    .Y(_07833_));
 sky130_fd_sc_hd__nand2_1 _14663_ (.A(_07409_),
    .B(_07833_),
    .Y(_07834_));
 sky130_fd_sc_hd__or2_1 _14664_ (.A(_07409_),
    .B(_07833_),
    .X(_07835_));
 sky130_fd_sc_hd__and2_1 _14665_ (.A(_07834_),
    .B(_07835_),
    .X(_07836_));
 sky130_fd_sc_hd__inv_2 _14666_ (.A(_07836_),
    .Y(_07837_));
 sky130_fd_sc_hd__inv_2 _14667_ (.A(_07471_),
    .Y(_07838_));
 sky130_fd_sc_hd__o21a_1 _14668_ (.A1(_07470_),
    .A2(_07527_),
    .B1(_07412_),
    .X(_07839_));
 sky130_fd_sc_hd__inv_2 _14669_ (.A(_07839_),
    .Y(_07840_));
 sky130_fd_sc_hd__o31a_2 _14670_ (.A1(_07838_),
    .A2(_07530_),
    .A3(_07802_),
    .B1(_07840_),
    .X(_07841_));
 sky130_fd_sc_hd__or3b_2 _14671_ (.A(_07404_),
    .B(_07406_),
    .C_N(_07832_),
    .X(_07842_));
 sky130_fd_sc_hd__a21oi_1 _14672_ (.A1(_06720_),
    .A2(_07829_),
    .B1(_07828_),
    .Y(_07843_));
 sky130_fd_sc_hd__clkinv_2 _14673_ (.A(_07402_),
    .Y(_07844_));
 sky130_fd_sc_hd__a2bb2o_1 _14674_ (.A1_N(_07830_),
    .A2_N(_07843_),
    .B1(_07831_),
    .B2(_07844_),
    .X(_07845_));
 sky130_fd_sc_hd__a21oi_2 _14675_ (.A1(_07830_),
    .A2(_07843_),
    .B1(_07845_),
    .Y(_07846_));
 sky130_fd_sc_hd__xnor2_2 _14676_ (.A(_07842_),
    .B(_07846_),
    .Y(_07847_));
 sky130_fd_sc_hd__inv_2 _14677_ (.A(_07847_),
    .Y(_07848_));
 sky130_fd_sc_hd__a21bo_1 _14678_ (.A1(_07842_),
    .A2(_07834_),
    .B1_N(_07846_),
    .X(_07849_));
 sky130_fd_sc_hd__o31ai_4 _14679_ (.A1(_07837_),
    .A2(_07841_),
    .A3(_07848_),
    .B1(_07849_),
    .Y(_07850_));
 sky130_fd_sc_hd__o21ba_1 _14680_ (.A1(_07206_),
    .A2(_07398_),
    .B1_N(_07337_),
    .X(_07851_));
 sky130_fd_sc_hd__and4b_1 _14681_ (.A_N(_07845_),
    .B(_07851_),
    .C(_07067_),
    .D(_07332_),
    .X(_07852_));
 sky130_fd_sc_hd__inv_2 _14682_ (.A(_07852_),
    .Y(_07853_));
 sky130_fd_sc_hd__xnor2_1 _14683_ (.A(_07850_),
    .B(_07853_),
    .Y(_07854_));
 sky130_fd_sc_hd__nand3_2 _14684_ (.A(_06613_),
    .B(_07850_),
    .C(_07853_),
    .Y(_07855_));
 sky130_fd_sc_hd__o21a_1 _14685_ (.A1(_07827_),
    .A2(_07854_),
    .B1(_07855_),
    .X(_07856_));
 sky130_fd_sc_hd__o21a_1 _14686_ (.A1(_07837_),
    .A2(_07841_),
    .B1(_07834_),
    .X(_07857_));
 sky130_fd_sc_hd__xnor2_2 _14687_ (.A(_07847_),
    .B(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__xnor2_1 _14688_ (.A(_07837_),
    .B(_07841_),
    .Y(_07859_));
 sky130_fd_sc_hd__nor2_1 _14689_ (.A(_06613_),
    .B(_07859_),
    .Y(_07860_));
 sky130_fd_sc_hd__a211o_1 _14690_ (.A1(_07827_),
    .A2(_07858_),
    .B1(_07860_),
    .C1(_07822_),
    .X(_07861_));
 sky130_fd_sc_hd__a21boi_2 _14691_ (.A1(_07822_),
    .A2(_07856_),
    .B1_N(_07861_),
    .Y(_07862_));
 sky130_fd_sc_hd__nand2_1 _14692_ (.A(_07067_),
    .B(_07826_),
    .Y(_07863_));
 sky130_fd_sc_hd__o211a_1 _14693_ (.A1(_07826_),
    .A2(_07862_),
    .B1(_07863_),
    .C1(_06568_),
    .X(_07864_));
 sky130_fd_sc_hd__o21ba_1 _14694_ (.A1(_06568_),
    .A2(_07825_),
    .B1_N(_07864_),
    .X(_07865_));
 sky130_fd_sc_hd__a21o_4 _14695_ (.A1(_06379_),
    .A2(_06505_),
    .B1(_06515_),
    .X(_07866_));
 sky130_fd_sc_hd__o21ai_4 _14696_ (.A1(_06470_),
    .A2(_07865_),
    .B1(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__and4b_2 _14697_ (.A_N(_04436_),
    .B(_04437_),
    .C(_04433_),
    .D(_06259_),
    .X(_07868_));
 sky130_fd_sc_hd__buf_4 _14698_ (.A(_07868_),
    .X(_07869_));
 sky130_fd_sc_hd__mux2_1 _14699_ (.A0(\rbzero.wall_tracer.stepDistY[-11] ),
    .A1(_07867_),
    .S(_07869_),
    .X(_07870_));
 sky130_fd_sc_hd__clkbuf_1 _14700_ (.A(_07870_),
    .X(_00391_));
 sky130_fd_sc_hd__and3_1 _14701_ (.A(_07806_),
    .B(_07850_),
    .C(_07853_),
    .X(_07871_));
 sky130_fd_sc_hd__xnor2_1 _14702_ (.A(_07850_),
    .B(_07852_),
    .Y(_07872_));
 sky130_fd_sc_hd__mux2_1 _14703_ (.A0(_07872_),
    .A1(_07858_),
    .S(_07806_),
    .X(_07873_));
 sky130_fd_sc_hd__mux2_1 _14704_ (.A0(_07871_),
    .A1(_07873_),
    .S(_06580_),
    .X(_07874_));
 sky130_fd_sc_hd__a21o_1 _14705_ (.A1(_06575_),
    .A2(_07874_),
    .B1(_06631_),
    .X(_07875_));
 sky130_fd_sc_hd__nor2_1 _14706_ (.A(_07806_),
    .B(_07859_),
    .Y(_07876_));
 sky130_fd_sc_hd__and2_1 _14707_ (.A(_07806_),
    .B(_07804_),
    .X(_07877_));
 sky130_fd_sc_hd__nor2_1 _14708_ (.A(_06613_),
    .B(_07809_),
    .Y(_07878_));
 sky130_fd_sc_hd__a21oi_1 _14709_ (.A1(_06613_),
    .A2(_07805_),
    .B1(_07878_),
    .Y(_07879_));
 sky130_fd_sc_hd__nand2_1 _14710_ (.A(_06580_),
    .B(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__o31a_1 _14711_ (.A1(_06580_),
    .A2(_07876_),
    .A3(_07877_),
    .B1(_07880_),
    .X(_07881_));
 sky130_fd_sc_hd__nor2_1 _14712_ (.A(_06579_),
    .B(_07819_),
    .Y(_07882_));
 sky130_fd_sc_hd__o21bai_1 _14713_ (.A1(_06613_),
    .A2(_07814_),
    .B1_N(_07882_),
    .Y(_07883_));
 sky130_fd_sc_hd__nor2_1 _14714_ (.A(_06579_),
    .B(_07808_),
    .Y(_07884_));
 sky130_fd_sc_hd__nor2_1 _14715_ (.A(_06613_),
    .B(_07817_),
    .Y(_07885_));
 sky130_fd_sc_hd__or2_1 _14716_ (.A(_07884_),
    .B(_07885_),
    .X(_07886_));
 sky130_fd_sc_hd__mux2_1 _14717_ (.A0(_07883_),
    .A1(_07886_),
    .S(_06584_),
    .X(_07887_));
 sky130_fd_sc_hd__or2_1 _14718_ (.A(_06595_),
    .B(_07887_),
    .X(_07888_));
 sky130_fd_sc_hd__o21a_1 _14719_ (.A1(_06575_),
    .A2(_07881_),
    .B1(_07888_),
    .X(_07889_));
 sky130_fd_sc_hd__or2_1 _14720_ (.A(_06568_),
    .B(_07889_),
    .X(_07890_));
 sky130_fd_sc_hd__clkbuf_4 _14721_ (.A(_06516_),
    .X(_07891_));
 sky130_fd_sc_hd__a31o_2 _14722_ (.A1(_06633_),
    .A2(_07875_),
    .A3(_07890_),
    .B1(_07891_),
    .X(_07892_));
 sky130_fd_sc_hd__mux2_1 _14723_ (.A0(\rbzero.wall_tracer.stepDistY[-10] ),
    .A1(_07892_),
    .S(_07869_),
    .X(_07893_));
 sky130_fd_sc_hd__clkbuf_1 _14724_ (.A(_07893_),
    .X(_00392_));
 sky130_fd_sc_hd__buf_2 _14725_ (.A(_06589_),
    .X(_07894_));
 sky130_fd_sc_hd__mux2_1 _14726_ (.A0(_07872_),
    .A1(_07858_),
    .S(_07827_),
    .X(_07895_));
 sky130_fd_sc_hd__or3b_1 _14727_ (.A(_06540_),
    .B(_06577_),
    .C_N(_07855_),
    .X(_07896_));
 sky130_fd_sc_hd__o211a_1 _14728_ (.A1(_07894_),
    .A2(_07895_),
    .B1(_07896_),
    .C1(_06619_),
    .X(_07897_));
 sky130_fd_sc_hd__nand2_1 _14729_ (.A(_07820_),
    .B(_07815_),
    .Y(_07898_));
 sky130_fd_sc_hd__xnor2_1 _14730_ (.A(_07836_),
    .B(_07841_),
    .Y(_07899_));
 sky130_fd_sc_hd__mux2_1 _14731_ (.A0(_07899_),
    .A1(_07804_),
    .S(_07827_),
    .X(_07900_));
 sky130_fd_sc_hd__a21o_1 _14732_ (.A1(_07806_),
    .A2(_07805_),
    .B1(_07810_),
    .X(_07901_));
 sky130_fd_sc_hd__mux2_1 _14733_ (.A0(_07900_),
    .A1(_07901_),
    .S(_06577_),
    .X(_07902_));
 sky130_fd_sc_hd__buf_2 _14734_ (.A(_06619_),
    .X(_07903_));
 sky130_fd_sc_hd__o21ai_1 _14735_ (.A1(_07827_),
    .A2(_07808_),
    .B1(_07818_),
    .Y(_07904_));
 sky130_fd_sc_hd__or2_1 _14736_ (.A(_06665_),
    .B(_07904_),
    .X(_07905_));
 sky130_fd_sc_hd__o221a_1 _14737_ (.A1(_06663_),
    .A2(_07898_),
    .B1(_07902_),
    .B2(_07903_),
    .C1(_07905_),
    .X(_07906_));
 sky130_fd_sc_hd__a221o_2 _14738_ (.A1(_06525_),
    .A2(_07897_),
    .B1(_07906_),
    .B2(_06670_),
    .C1(_07891_),
    .X(_07907_));
 sky130_fd_sc_hd__mux2_1 _14739_ (.A0(\rbzero.wall_tracer.stepDistY[-9] ),
    .A1(_07907_),
    .S(_07869_),
    .X(_07908_));
 sky130_fd_sc_hd__clkbuf_1 _14740_ (.A(_07908_),
    .X(_00393_));
 sky130_fd_sc_hd__a21oi_1 _14741_ (.A1(_07806_),
    .A2(_07858_),
    .B1(_07876_),
    .Y(_07909_));
 sky130_fd_sc_hd__and2_1 _14742_ (.A(_07827_),
    .B(_07805_),
    .X(_07910_));
 sky130_fd_sc_hd__a21oi_1 _14743_ (.A1(_07806_),
    .A2(_07804_),
    .B1(_07910_),
    .Y(_07911_));
 sky130_fd_sc_hd__and2_1 _14744_ (.A(_06577_),
    .B(_07911_),
    .X(_07912_));
 sky130_fd_sc_hd__a211o_1 _14745_ (.A1(_07894_),
    .A2(_07909_),
    .B1(_07912_),
    .C1(_07903_),
    .X(_07913_));
 sky130_fd_sc_hd__nor2_1 _14746_ (.A(_07878_),
    .B(_07884_),
    .Y(_07914_));
 sky130_fd_sc_hd__nor2_1 _14747_ (.A(_07885_),
    .B(_07882_),
    .Y(_07915_));
 sky130_fd_sc_hd__o221a_1 _14748_ (.A1(_06665_),
    .A2(_07914_),
    .B1(_07915_),
    .B2(_06663_),
    .C1(_06602_),
    .X(_07916_));
 sky130_fd_sc_hd__a21o_1 _14749_ (.A1(_07827_),
    .A2(_07872_),
    .B1(_07871_),
    .X(_07917_));
 sky130_fd_sc_hd__a21oi_1 _14750_ (.A1(_06598_),
    .A2(_07917_),
    .B1(_06602_),
    .Y(_07918_));
 sky130_fd_sc_hd__a211o_1 _14751_ (.A1(_07913_),
    .A2(_07916_),
    .B1(_07918_),
    .C1(_06470_),
    .X(_07919_));
 sky130_fd_sc_hd__nand2_1 _14752_ (.A(_07822_),
    .B(_07883_),
    .Y(_07920_));
 sky130_fd_sc_hd__nor2_1 _14753_ (.A(_06574_),
    .B(_07920_),
    .Y(_07921_));
 sky130_fd_sc_hd__a21oi_1 _14754_ (.A1(_06655_),
    .A2(_07921_),
    .B1(_07891_),
    .Y(_07922_));
 sky130_fd_sc_hd__nand2_2 _14755_ (.A(_07919_),
    .B(_07922_),
    .Y(_07923_));
 sky130_fd_sc_hd__mux2_1 _14756_ (.A0(\rbzero.wall_tracer.stepDistY[-8] ),
    .A1(_07923_),
    .S(_07869_),
    .X(_07924_));
 sky130_fd_sc_hd__clkbuf_1 _14757_ (.A(_07924_),
    .X(_00394_));
 sky130_fd_sc_hd__xnor2_1 _14758_ (.A(_07848_),
    .B(_07857_),
    .Y(_07925_));
 sky130_fd_sc_hd__mux2_1 _14759_ (.A0(_07854_),
    .A1(_07925_),
    .S(_07827_),
    .X(_07926_));
 sky130_fd_sc_hd__nor2_1 _14760_ (.A(_07894_),
    .B(_07900_),
    .Y(_07927_));
 sky130_fd_sc_hd__a211o_1 _14761_ (.A1(_07894_),
    .A2(_07926_),
    .B1(_07927_),
    .C1(_07903_),
    .X(_07928_));
 sky130_fd_sc_hd__mux2_1 _14762_ (.A0(_07904_),
    .A1(_07901_),
    .S(_07894_),
    .X(_07929_));
 sky130_fd_sc_hd__a21oi_1 _14763_ (.A1(_07903_),
    .A2(_07929_),
    .B1(_06669_),
    .Y(_07930_));
 sky130_fd_sc_hd__a21o_1 _14764_ (.A1(_07067_),
    .A2(_07855_),
    .B1(_06663_),
    .X(_07931_));
 sky130_fd_sc_hd__a21o_1 _14765_ (.A1(_06669_),
    .A2(_07931_),
    .B1(_06470_),
    .X(_07932_));
 sky130_fd_sc_hd__a21o_1 _14766_ (.A1(_07928_),
    .A2(_07930_),
    .B1(_07932_),
    .X(_07933_));
 sky130_fd_sc_hd__a31oi_2 _14767_ (.A1(_06470_),
    .A2(_07826_),
    .A3(_07823_),
    .B1(_07891_),
    .Y(_07934_));
 sky130_fd_sc_hd__nand2_2 _14768_ (.A(_07933_),
    .B(_07934_),
    .Y(_07935_));
 sky130_fd_sc_hd__mux2_1 _14769_ (.A0(\rbzero.wall_tracer.stepDistY[-7] ),
    .A1(_07935_),
    .S(_07869_),
    .X(_07936_));
 sky130_fd_sc_hd__clkbuf_1 _14770_ (.A(_07936_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _14771_ (.A0(_07914_),
    .A1(_07911_),
    .S(_07894_),
    .X(_07937_));
 sky130_fd_sc_hd__a211o_1 _14772_ (.A1(_07827_),
    .A2(_07872_),
    .B1(_07871_),
    .C1(_06577_),
    .X(_07938_));
 sky130_fd_sc_hd__a211o_1 _14773_ (.A1(_07806_),
    .A2(_07858_),
    .B1(_07876_),
    .C1(_06589_),
    .X(_07939_));
 sky130_fd_sc_hd__a21oi_1 _14774_ (.A1(_07938_),
    .A2(_07939_),
    .B1(_07903_),
    .Y(_07940_));
 sky130_fd_sc_hd__nand2_1 _14775_ (.A(_06633_),
    .B(_06602_),
    .Y(_07941_));
 sky130_fd_sc_hd__a211oi_2 _14776_ (.A1(_07903_),
    .A2(_07937_),
    .B1(_07940_),
    .C1(_07941_),
    .Y(_07942_));
 sky130_fd_sc_hd__and3_1 _14777_ (.A(_06655_),
    .B(_07826_),
    .C(_07887_),
    .X(_07943_));
 sky130_fd_sc_hd__or3_2 _14778_ (.A(_07891_),
    .B(_07942_),
    .C(_07943_),
    .X(_07944_));
 sky130_fd_sc_hd__mux2_1 _14779_ (.A0(\rbzero.wall_tracer.stepDistY[-6] ),
    .A1(_07944_),
    .S(_07869_),
    .X(_07945_));
 sky130_fd_sc_hd__clkbuf_1 _14780_ (.A(_07945_),
    .X(_00396_));
 sky130_fd_sc_hd__or2_1 _14781_ (.A(_06577_),
    .B(_07855_),
    .X(_07946_));
 sky130_fd_sc_hd__o211a_1 _14782_ (.A1(_07894_),
    .A2(_07926_),
    .B1(_07946_),
    .C1(_06641_),
    .X(_07947_));
 sky130_fd_sc_hd__o21ai_1 _14783_ (.A1(_06641_),
    .A2(_07902_),
    .B1(_06670_),
    .Y(_07948_));
 sky130_fd_sc_hd__nor2_1 _14784_ (.A(_07822_),
    .B(_07821_),
    .Y(_07949_));
 sky130_fd_sc_hd__a21o_1 _14785_ (.A1(_07822_),
    .A2(_07811_),
    .B1(_07949_),
    .X(_07950_));
 sky130_fd_sc_hd__or2_1 _14786_ (.A(_06580_),
    .B(_07815_),
    .X(_07951_));
 sky130_fd_sc_hd__mux2_1 _14787_ (.A0(_07950_),
    .A1(_07951_),
    .S(_06574_),
    .X(_07952_));
 sky130_fd_sc_hd__o21a_1 _14788_ (.A1(_06581_),
    .A2(_07952_),
    .B1(_07866_),
    .X(_07953_));
 sky130_fd_sc_hd__o21ai_4 _14789_ (.A1(_07947_),
    .A2(_07948_),
    .B1(_07953_),
    .Y(_07954_));
 sky130_fd_sc_hd__mux2_1 _14790_ (.A0(\rbzero.wall_tracer.stepDistY[-5] ),
    .A1(_07954_),
    .S(_07869_),
    .X(_07955_));
 sky130_fd_sc_hd__clkbuf_1 _14791_ (.A(_07955_),
    .X(_00397_));
 sky130_fd_sc_hd__a21o_1 _14792_ (.A1(_07894_),
    .A2(_07909_),
    .B1(_07912_),
    .X(_07956_));
 sky130_fd_sc_hd__a21oi_1 _14793_ (.A1(_06577_),
    .A2(_07917_),
    .B1(_07903_),
    .Y(_07957_));
 sky130_fd_sc_hd__a211o_1 _14794_ (.A1(_07903_),
    .A2(_07956_),
    .B1(_07957_),
    .C1(_07941_),
    .X(_07958_));
 sky130_fd_sc_hd__nor2_1 _14795_ (.A(_07822_),
    .B(_07886_),
    .Y(_07959_));
 sky130_fd_sc_hd__and2_1 _14796_ (.A(_07822_),
    .B(_07879_),
    .X(_07960_));
 sky130_fd_sc_hd__or2_1 _14797_ (.A(_07826_),
    .B(_07920_),
    .X(_07961_));
 sky130_fd_sc_hd__o31a_1 _14798_ (.A1(_06574_),
    .A2(_07959_),
    .A3(_07960_),
    .B1(_07961_),
    .X(_07962_));
 sky130_fd_sc_hd__or2_1 _14799_ (.A(_06581_),
    .B(_07962_),
    .X(_07963_));
 sky130_fd_sc_hd__nand3_2 _14800_ (.A(_07866_),
    .B(_07958_),
    .C(_07963_),
    .Y(_07964_));
 sky130_fd_sc_hd__mux2_1 _14801_ (.A0(\rbzero.wall_tracer.stepDistY[-4] ),
    .A1(_07964_),
    .S(_07869_),
    .X(_07965_));
 sky130_fd_sc_hd__clkbuf_1 _14802_ (.A(_07965_),
    .X(_00398_));
 sky130_fd_sc_hd__a21o_1 _14803_ (.A1(_07894_),
    .A2(_07926_),
    .B1(_07927_),
    .X(_07966_));
 sky130_fd_sc_hd__a21oi_1 _14804_ (.A1(_07067_),
    .A2(_07855_),
    .B1(_07894_),
    .Y(_07967_));
 sky130_fd_sc_hd__nor2_1 _14805_ (.A(_07903_),
    .B(_07967_),
    .Y(_07968_));
 sky130_fd_sc_hd__a211oi_2 _14806_ (.A1(_07903_),
    .A2(_07966_),
    .B1(_07968_),
    .C1(_07941_),
    .Y(_07969_));
 sky130_fd_sc_hd__o21ai_1 _14807_ (.A1(_06581_),
    .A2(_07825_),
    .B1(_07866_),
    .Y(_07970_));
 sky130_fd_sc_hd__or2_2 _14808_ (.A(_07969_),
    .B(_07970_),
    .X(_07971_));
 sky130_fd_sc_hd__mux2_1 _14809_ (.A0(\rbzero.wall_tracer.stepDistY[-3] ),
    .A1(_07971_),
    .S(_07869_),
    .X(_07972_));
 sky130_fd_sc_hd__clkbuf_1 _14810_ (.A(_07972_),
    .X(_00399_));
 sky130_fd_sc_hd__and3_1 _14811_ (.A(_06619_),
    .B(_07938_),
    .C(_07939_),
    .X(_07973_));
 sky130_fd_sc_hd__o211a_1 _14812_ (.A1(_06574_),
    .A2(_07881_),
    .B1(_07888_),
    .C1(_06655_),
    .X(_07974_));
 sky130_fd_sc_hd__a211o_4 _14813_ (.A1(_06670_),
    .A2(_07973_),
    .B1(_07974_),
    .C1(_06516_),
    .X(_07975_));
 sky130_fd_sc_hd__mux2_1 _14814_ (.A0(\rbzero.wall_tracer.stepDistY[-2] ),
    .A1(_07975_),
    .S(_07869_),
    .X(_07976_));
 sky130_fd_sc_hd__clkbuf_1 _14815_ (.A(_07976_),
    .X(_00400_));
 sky130_fd_sc_hd__or2_1 _14816_ (.A(_07822_),
    .B(_07807_),
    .X(_07977_));
 sky130_fd_sc_hd__a211o_1 _14817_ (.A1(_07827_),
    .A2(_07858_),
    .B1(_07860_),
    .C1(_06580_),
    .X(_07978_));
 sky130_fd_sc_hd__nor2_1 _14818_ (.A(_06595_),
    .B(_07950_),
    .Y(_07979_));
 sky130_fd_sc_hd__a311o_1 _14819_ (.A1(_06595_),
    .A2(_07977_),
    .A3(_07978_),
    .B1(_07979_),
    .C1(_06631_),
    .X(_07980_));
 sky130_fd_sc_hd__a22oi_4 _14820_ (.A1(_06602_),
    .A2(_07897_),
    .B1(_07980_),
    .B2(_06655_),
    .Y(_07981_));
 sky130_fd_sc_hd__nand2_4 _14821_ (.A(_07866_),
    .B(_07981_),
    .Y(_07982_));
 sky130_fd_sc_hd__buf_4 _14822_ (.A(_07868_),
    .X(_07983_));
 sky130_fd_sc_hd__mux2_1 _14823_ (.A0(\rbzero.wall_tracer.stepDistY[-1] ),
    .A1(_07982_),
    .S(_07983_),
    .X(_07984_));
 sky130_fd_sc_hd__clkbuf_1 _14824_ (.A(_07984_),
    .X(_00401_));
 sky130_fd_sc_hd__or2_1 _14825_ (.A(_07876_),
    .B(_07877_),
    .X(_07985_));
 sky130_fd_sc_hd__mux2_1 _14826_ (.A0(_07873_),
    .A1(_07985_),
    .S(_06580_),
    .X(_07986_));
 sky130_fd_sc_hd__or3_1 _14827_ (.A(_06595_),
    .B(_07959_),
    .C(_07960_),
    .X(_07987_));
 sky130_fd_sc_hd__a21bo_1 _14828_ (.A1(_07826_),
    .A2(_07986_),
    .B1_N(_07987_),
    .X(_07988_));
 sky130_fd_sc_hd__nor2_2 _14829_ (.A(_06515_),
    .B(_06498_),
    .Y(_07989_));
 sky130_fd_sc_hd__and2_1 _14830_ (.A(_07989_),
    .B(_07921_),
    .X(_07990_));
 sky130_fd_sc_hd__a31o_1 _14831_ (.A1(_06602_),
    .A2(_06598_),
    .A3(_07917_),
    .B1(_06516_),
    .X(_07991_));
 sky130_fd_sc_hd__a211o_4 _14832_ (.A1(_06655_),
    .A2(_07988_),
    .B1(_07990_),
    .C1(_07991_),
    .X(_07992_));
 sky130_fd_sc_hd__mux2_1 _14833_ (.A0(\rbzero.wall_tracer.stepDistY[0] ),
    .A1(_07992_),
    .S(_07983_),
    .X(_07993_));
 sky130_fd_sc_hd__clkbuf_1 _14834_ (.A(_07993_),
    .X(_00402_));
 sky130_fd_sc_hd__nand2_1 _14835_ (.A(_06575_),
    .B(_07813_),
    .Y(_07994_));
 sky130_fd_sc_hd__o21ai_2 _14836_ (.A1(_06575_),
    .A2(_07862_),
    .B1(_07994_),
    .Y(_07995_));
 sky130_fd_sc_hd__o221ai_4 _14837_ (.A1(_06669_),
    .A2(_07931_),
    .B1(_07995_),
    .B2(_06581_),
    .C1(_07866_),
    .Y(_07996_));
 sky130_fd_sc_hd__mux2_1 _14838_ (.A0(\rbzero.wall_tracer.stepDistY[1] ),
    .A1(_07996_),
    .S(_07983_),
    .X(_07997_));
 sky130_fd_sc_hd__clkbuf_1 _14839_ (.A(_07997_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _14840_ (.A0(_07874_),
    .A1(_07881_),
    .S(_06575_),
    .X(_07998_));
 sky130_fd_sc_hd__a31o_1 _14841_ (.A1(_07826_),
    .A2(_07989_),
    .A3(_07887_),
    .B1(_06516_),
    .X(_07999_));
 sky130_fd_sc_hd__a21o_4 _14842_ (.A1(_06655_),
    .A2(_07998_),
    .B1(_07999_),
    .X(_08000_));
 sky130_fd_sc_hd__mux2_1 _14843_ (.A0(\rbzero.wall_tracer.stepDistY[2] ),
    .A1(_08000_),
    .S(_07983_),
    .X(_08001_));
 sky130_fd_sc_hd__clkbuf_1 _14844_ (.A(_08001_),
    .X(_00404_));
 sky130_fd_sc_hd__nand2_1 _14845_ (.A(_06631_),
    .B(_07952_),
    .Y(_08002_));
 sky130_fd_sc_hd__nor2_1 _14846_ (.A(_07822_),
    .B(_07856_),
    .Y(_08003_));
 sky130_fd_sc_hd__a31o_1 _14847_ (.A1(_06574_),
    .A2(_07977_),
    .A3(_07978_),
    .B1(_06631_),
    .X(_08004_));
 sky130_fd_sc_hd__a21o_1 _14848_ (.A1(_07826_),
    .A2(_08003_),
    .B1(_08004_),
    .X(_08005_));
 sky130_fd_sc_hd__a31o_2 _14849_ (.A1(_06470_),
    .A2(_08002_),
    .A3(_08005_),
    .B1(_06516_),
    .X(_08006_));
 sky130_fd_sc_hd__mux2_1 _14850_ (.A0(\rbzero.wall_tracer.stepDistY[3] ),
    .A1(_08006_),
    .S(_07983_),
    .X(_08007_));
 sky130_fd_sc_hd__clkbuf_1 _14851_ (.A(_08007_),
    .X(_00405_));
 sky130_fd_sc_hd__a31o_1 _14852_ (.A1(_06577_),
    .A2(_07826_),
    .A3(_07871_),
    .B1(_06631_),
    .X(_08008_));
 sky130_fd_sc_hd__a21o_1 _14853_ (.A1(_06575_),
    .A2(_07986_),
    .B1(_08008_),
    .X(_08009_));
 sky130_fd_sc_hd__nand2_1 _14854_ (.A(_06631_),
    .B(_07962_),
    .Y(_08010_));
 sky130_fd_sc_hd__a31o_1 _14855_ (.A1(_06470_),
    .A2(_08009_),
    .A3(_08010_),
    .B1(_07891_),
    .X(_08011_));
 sky130_fd_sc_hd__buf_2 _14856_ (.A(_08011_),
    .X(_08012_));
 sky130_fd_sc_hd__mux2_1 _14857_ (.A0(\rbzero.wall_tracer.stepDistY[4] ),
    .A1(_08012_),
    .S(_07983_),
    .X(_08013_));
 sky130_fd_sc_hd__clkbuf_1 _14858_ (.A(_08013_),
    .X(_00406_));
 sky130_fd_sc_hd__o21ai_1 _14859_ (.A1(_06600_),
    .A2(_07825_),
    .B1(_07866_),
    .Y(_08014_));
 sky130_fd_sc_hd__a31o_1 _14860_ (.A1(_06470_),
    .A2(_06575_),
    .A3(_07862_),
    .B1(_08014_),
    .X(_08015_));
 sky130_fd_sc_hd__mux2_1 _14861_ (.A0(\rbzero.wall_tracer.stepDistY[5] ),
    .A1(_08015_),
    .S(_07983_),
    .X(_08016_));
 sky130_fd_sc_hd__clkbuf_1 _14862_ (.A(_08016_),
    .X(_00407_));
 sky130_fd_sc_hd__a21o_1 _14863_ (.A1(_07989_),
    .A2(_07889_),
    .B1(_06516_),
    .X(_08017_));
 sky130_fd_sc_hd__a31o_1 _14864_ (.A1(_06470_),
    .A2(_06575_),
    .A3(_07874_),
    .B1(_08017_),
    .X(_08018_));
 sky130_fd_sc_hd__mux2_1 _14865_ (.A0(\rbzero.wall_tracer.stepDistY[6] ),
    .A1(_08018_),
    .S(_07983_),
    .X(_08019_));
 sky130_fd_sc_hd__clkbuf_1 _14866_ (.A(_08019_),
    .X(_00408_));
 sky130_fd_sc_hd__a31o_1 _14867_ (.A1(_07826_),
    .A2(_07977_),
    .A3(_07978_),
    .B1(_07979_),
    .X(_08020_));
 sky130_fd_sc_hd__or2_1 _14868_ (.A(_06568_),
    .B(_08020_),
    .X(_08021_));
 sky130_fd_sc_hd__a31o_1 _14869_ (.A1(_06470_),
    .A2(_06575_),
    .A3(_08003_),
    .B1(_07989_),
    .X(_08022_));
 sky130_fd_sc_hd__a21o_1 _14870_ (.A1(_08021_),
    .A2(_08022_),
    .B1(_07891_),
    .X(_08023_));
 sky130_fd_sc_hd__mux2_1 _14871_ (.A0(\rbzero.wall_tracer.stepDistY[7] ),
    .A1(_08023_),
    .S(_07983_),
    .X(_08024_));
 sky130_fd_sc_hd__clkbuf_1 _14872_ (.A(_08024_),
    .X(_00409_));
 sky130_fd_sc_hd__a31o_1 _14873_ (.A1(_06470_),
    .A2(_06598_),
    .A3(_07871_),
    .B1(_07989_),
    .X(_08025_));
 sky130_fd_sc_hd__o21a_1 _14874_ (.A1(_06568_),
    .A2(_07988_),
    .B1(_08025_),
    .X(_08026_));
 sky130_fd_sc_hd__or2_1 _14875_ (.A(_07891_),
    .B(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__mux2_1 _14876_ (.A0(\rbzero.wall_tracer.stepDistY[8] ),
    .A1(_08027_),
    .S(_07983_),
    .X(_08028_));
 sky130_fd_sc_hd__clkbuf_1 _14877_ (.A(_08028_),
    .X(_00410_));
 sky130_fd_sc_hd__o21ai_2 _14878_ (.A1(_06600_),
    .A2(_07995_),
    .B1(_07866_),
    .Y(_08029_));
 sky130_fd_sc_hd__mux2_1 _14879_ (.A0(\rbzero.wall_tracer.stepDistY[9] ),
    .A1(_08029_),
    .S(_07868_),
    .X(_08030_));
 sky130_fd_sc_hd__clkbuf_1 _14880_ (.A(_08030_),
    .X(_00411_));
 sky130_fd_sc_hd__and4bb_1 _14881_ (.A_N(_07891_),
    .B_N(_06541_),
    .C(_06631_),
    .D(_07998_),
    .X(_08031_));
 sky130_fd_sc_hd__mux2_1 _14882_ (.A0(\rbzero.wall_tracer.stepDistY[10] ),
    .A1(_08031_),
    .S(_07868_),
    .X(_08032_));
 sky130_fd_sc_hd__clkbuf_1 _14883_ (.A(_08032_),
    .X(_00412_));
 sky130_fd_sc_hd__nand2_4 _14884_ (.A(_06160_),
    .B(_06257_),
    .Y(_08033_));
 sky130_fd_sc_hd__or2_1 _14885_ (.A(_06103_),
    .B(_08033_),
    .X(_08034_));
 sky130_fd_sc_hd__clkbuf_4 _14886_ (.A(_08034_),
    .X(_08035_));
 sky130_fd_sc_hd__clkbuf_4 _14887_ (.A(_08035_),
    .X(_08036_));
 sky130_fd_sc_hd__buf_4 _14888_ (.A(_06217_),
    .X(_08037_));
 sky130_fd_sc_hd__mux2_1 _14889_ (.A0(\rbzero.wall_tracer.trackDistY[-11] ),
    .A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .S(_08037_),
    .X(_08038_));
 sky130_fd_sc_hd__inv_2 _14890_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .Y(_08039_));
 sky130_fd_sc_hd__nand2_1 _14891_ (.A(_08039_),
    .B(_08035_),
    .Y(_08040_));
 sky130_fd_sc_hd__buf_4 _14892_ (.A(_04442_),
    .X(_01633_));
 sky130_fd_sc_hd__o211a_1 _14893_ (.A1(_08036_),
    .A2(_08038_),
    .B1(_08040_),
    .C1(_01633_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _14894_ (.A0(\rbzero.wall_tracer.trackDistY[-10] ),
    .A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .S(_08037_),
    .X(_08041_));
 sky130_fd_sc_hd__inv_2 _14895_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .Y(_08042_));
 sky130_fd_sc_hd__nand2_1 _14896_ (.A(_08042_),
    .B(_08035_),
    .Y(_08043_));
 sky130_fd_sc_hd__o211a_1 _14897_ (.A1(_08036_),
    .A2(_08041_),
    .B1(_08043_),
    .C1(_01633_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _14898_ (.A0(\rbzero.wall_tracer.trackDistY[-9] ),
    .A1(\rbzero.wall_tracer.trackDistX[-9] ),
    .S(_08037_),
    .X(_08044_));
 sky130_fd_sc_hd__nor2_1 _14899_ (.A(_06103_),
    .B(_08033_),
    .Y(_08045_));
 sky130_fd_sc_hd__buf_2 _14900_ (.A(_08045_),
    .X(_08046_));
 sky130_fd_sc_hd__buf_2 _14901_ (.A(_08046_),
    .X(_08047_));
 sky130_fd_sc_hd__or2_1 _14902_ (.A(\rbzero.wall_tracer.visualWallDist[-9] ),
    .B(_08047_),
    .X(_08048_));
 sky130_fd_sc_hd__o211a_1 _14903_ (.A1(_08036_),
    .A2(_08044_),
    .B1(_08048_),
    .C1(_01633_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _14904_ (.A0(\rbzero.wall_tracer.trackDistY[-8] ),
    .A1(\rbzero.wall_tracer.trackDistX[-8] ),
    .S(_08037_),
    .X(_08049_));
 sky130_fd_sc_hd__or2_1 _14905_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(_08047_),
    .X(_08050_));
 sky130_fd_sc_hd__o211a_1 _14906_ (.A1(_08036_),
    .A2(_08049_),
    .B1(_08050_),
    .C1(_01633_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _14907_ (.A0(\rbzero.wall_tracer.trackDistY[-7] ),
    .A1(\rbzero.wall_tracer.trackDistX[-7] ),
    .S(_08037_),
    .X(_08051_));
 sky130_fd_sc_hd__or2_1 _14908_ (.A(\rbzero.wall_tracer.visualWallDist[-7] ),
    .B(_08047_),
    .X(_08052_));
 sky130_fd_sc_hd__o211a_1 _14909_ (.A1(_08036_),
    .A2(_08051_),
    .B1(_08052_),
    .C1(_01633_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _14910_ (.A0(\rbzero.wall_tracer.trackDistY[-6] ),
    .A1(\rbzero.wall_tracer.trackDistX[-6] ),
    .S(_08037_),
    .X(_08053_));
 sky130_fd_sc_hd__or2_1 _14911_ (.A(\rbzero.wall_tracer.visualWallDist[-6] ),
    .B(_08047_),
    .X(_08054_));
 sky130_fd_sc_hd__o211a_1 _14912_ (.A1(_08036_),
    .A2(_08053_),
    .B1(_08054_),
    .C1(_01633_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _14913_ (.A0(\rbzero.wall_tracer.trackDistY[-5] ),
    .A1(\rbzero.wall_tracer.trackDistX[-5] ),
    .S(_08037_),
    .X(_08055_));
 sky130_fd_sc_hd__or2_1 _14914_ (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .B(_08047_),
    .X(_08056_));
 sky130_fd_sc_hd__o211a_1 _14915_ (.A1(_08036_),
    .A2(_08055_),
    .B1(_08056_),
    .C1(_01633_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _14916_ (.A0(\rbzero.wall_tracer.trackDistY[-4] ),
    .A1(\rbzero.wall_tracer.trackDistX[-4] ),
    .S(_08037_),
    .X(_08057_));
 sky130_fd_sc_hd__or2_1 _14917_ (.A(\rbzero.wall_tracer.visualWallDist[-4] ),
    .B(_08047_),
    .X(_08058_));
 sky130_fd_sc_hd__o211a_1 _14918_ (.A1(_08036_),
    .A2(_08057_),
    .B1(_08058_),
    .C1(_01633_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _14919_ (.A0(\rbzero.wall_tracer.trackDistY[-3] ),
    .A1(\rbzero.wall_tracer.trackDistX[-3] ),
    .S(_08037_),
    .X(_08059_));
 sky130_fd_sc_hd__or2_1 _14920_ (.A(\rbzero.wall_tracer.visualWallDist[-3] ),
    .B(_08047_),
    .X(_08060_));
 sky130_fd_sc_hd__buf_2 _14921_ (.A(_04442_),
    .X(_08061_));
 sky130_fd_sc_hd__o211a_1 _14922_ (.A1(_08036_),
    .A2(_08059_),
    .B1(_08060_),
    .C1(_08061_),
    .X(_00421_));
 sky130_fd_sc_hd__clkbuf_4 _14923_ (.A(_06217_),
    .X(_08062_));
 sky130_fd_sc_hd__mux2_1 _14924_ (.A0(\rbzero.wall_tracer.trackDistY[-2] ),
    .A1(\rbzero.wall_tracer.trackDistX[-2] ),
    .S(_08062_),
    .X(_08063_));
 sky130_fd_sc_hd__or2_1 _14925_ (.A(\rbzero.wall_tracer.visualWallDist[-2] ),
    .B(_08047_),
    .X(_08064_));
 sky130_fd_sc_hd__o211a_1 _14926_ (.A1(_08036_),
    .A2(_08063_),
    .B1(_08064_),
    .C1(_08061_),
    .X(_00422_));
 sky130_fd_sc_hd__buf_2 _14927_ (.A(_08035_),
    .X(_08065_));
 sky130_fd_sc_hd__mux2_1 _14928_ (.A0(\rbzero.wall_tracer.trackDistY[-1] ),
    .A1(\rbzero.wall_tracer.trackDistX[-1] ),
    .S(_08062_),
    .X(_08066_));
 sky130_fd_sc_hd__or2_1 _14929_ (.A(\rbzero.wall_tracer.visualWallDist[-1] ),
    .B(_08046_),
    .X(_08067_));
 sky130_fd_sc_hd__o211a_1 _14930_ (.A1(_08065_),
    .A2(_08066_),
    .B1(_08067_),
    .C1(_08061_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _14931_ (.A0(\rbzero.wall_tracer.trackDistY[0] ),
    .A1(\rbzero.wall_tracer.trackDistX[0] ),
    .S(_08062_),
    .X(_08068_));
 sky130_fd_sc_hd__inv_2 _14932_ (.A(\rbzero.wall_tracer.visualWallDist[0] ),
    .Y(_08069_));
 sky130_fd_sc_hd__nand2_1 _14933_ (.A(_08069_),
    .B(_08035_),
    .Y(_08070_));
 sky130_fd_sc_hd__o211a_1 _14934_ (.A1(_08065_),
    .A2(_08068_),
    .B1(_08070_),
    .C1(_08061_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _14935_ (.A0(\rbzero.wall_tracer.trackDistY[1] ),
    .A1(\rbzero.wall_tracer.trackDistX[1] ),
    .S(_08062_),
    .X(_08071_));
 sky130_fd_sc_hd__or2_1 _14936_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08046_),
    .X(_08072_));
 sky130_fd_sc_hd__o211a_1 _14937_ (.A1(_08065_),
    .A2(_08071_),
    .B1(_08072_),
    .C1(_08061_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _14938_ (.A0(\rbzero.wall_tracer.trackDistY[2] ),
    .A1(\rbzero.wall_tracer.trackDistX[2] ),
    .S(_08062_),
    .X(_08073_));
 sky130_fd_sc_hd__or2_1 _14939_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08046_),
    .X(_08074_));
 sky130_fd_sc_hd__o211a_1 _14940_ (.A1(_08065_),
    .A2(_08073_),
    .B1(_08074_),
    .C1(_08061_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _14941_ (.A0(\rbzero.wall_tracer.trackDistY[3] ),
    .A1(\rbzero.wall_tracer.trackDistX[3] ),
    .S(_08062_),
    .X(_08075_));
 sky130_fd_sc_hd__or2_1 _14942_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08046_),
    .X(_08076_));
 sky130_fd_sc_hd__o211a_1 _14943_ (.A1(_08065_),
    .A2(_08075_),
    .B1(_08076_),
    .C1(_08061_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _14944_ (.A0(\rbzero.wall_tracer.trackDistY[4] ),
    .A1(\rbzero.wall_tracer.trackDistX[4] ),
    .S(_08062_),
    .X(_08077_));
 sky130_fd_sc_hd__or2_1 _14945_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08046_),
    .X(_08078_));
 sky130_fd_sc_hd__o211a_1 _14946_ (.A1(_08065_),
    .A2(_08077_),
    .B1(_08078_),
    .C1(_08061_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _14947_ (.A0(\rbzero.wall_tracer.trackDistY[5] ),
    .A1(\rbzero.wall_tracer.trackDistX[5] ),
    .S(_08062_),
    .X(_08079_));
 sky130_fd_sc_hd__or2_1 _14948_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08046_),
    .X(_08080_));
 sky130_fd_sc_hd__o211a_1 _14949_ (.A1(_08065_),
    .A2(_08079_),
    .B1(_08080_),
    .C1(_08061_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _14950_ (.A0(\rbzero.wall_tracer.trackDistY[6] ),
    .A1(\rbzero.wall_tracer.trackDistX[6] ),
    .S(_08062_),
    .X(_08081_));
 sky130_fd_sc_hd__or2_1 _14951_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08046_),
    .X(_08082_));
 sky130_fd_sc_hd__o211a_1 _14952_ (.A1(_08065_),
    .A2(_08081_),
    .B1(_08082_),
    .C1(_08061_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _14953_ (.A0(\rbzero.wall_tracer.trackDistY[7] ),
    .A1(\rbzero.wall_tracer.trackDistX[7] ),
    .S(_08062_),
    .X(_08083_));
 sky130_fd_sc_hd__or2_1 _14954_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_08046_),
    .X(_08084_));
 sky130_fd_sc_hd__clkbuf_8 _14955_ (.A(_04442_),
    .X(_08085_));
 sky130_fd_sc_hd__o211a_1 _14956_ (.A1(_08065_),
    .A2(_08083_),
    .B1(_08084_),
    .C1(_08085_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _14957_ (.A0(\rbzero.wall_tracer.trackDistY[8] ),
    .A1(\rbzero.wall_tracer.trackDistX[8] ),
    .S(_06217_),
    .X(_08086_));
 sky130_fd_sc_hd__or2_1 _14958_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_08046_),
    .X(_08087_));
 sky130_fd_sc_hd__o211a_1 _14959_ (.A1(_08065_),
    .A2(_08086_),
    .B1(_08087_),
    .C1(_08085_),
    .X(_00432_));
 sky130_fd_sc_hd__nor3b_1 _14960_ (.A(_06215_),
    .B(_06216_),
    .C_N(\rbzero.wall_tracer.trackDistY[9] ),
    .Y(_08088_));
 sky130_fd_sc_hd__a211o_1 _14961_ (.A1(\rbzero.wall_tracer.trackDistX[9] ),
    .A2(_08037_),
    .B1(_08035_),
    .C1(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__o211a_1 _14962_ (.A1(\rbzero.wall_tracer.visualWallDist[9] ),
    .A2(_08047_),
    .B1(_08089_),
    .C1(_08085_),
    .X(_00433_));
 sky130_fd_sc_hd__a21o_1 _14963_ (.A1(\rbzero.wall_tracer.trackDistX[10] ),
    .A2(\rbzero.wall_tracer.trackDistY[10] ),
    .B1(_08035_),
    .X(_08090_));
 sky130_fd_sc_hd__o211a_1 _14964_ (.A1(\rbzero.wall_tracer.visualWallDist[10] ),
    .A2(_08047_),
    .B1(_08090_),
    .C1(_08085_),
    .X(_00434_));
 sky130_fd_sc_hd__and4b_2 _14965_ (.A_N(_04437_),
    .B(_04433_),
    .C(_04438_),
    .D(_04436_),
    .X(_08091_));
 sky130_fd_sc_hd__buf_4 _14966_ (.A(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__mux2_1 _14967_ (.A0(\rbzero.wall_tracer.stepDistX[-11] ),
    .A1(_07867_),
    .S(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__clkbuf_1 _14968_ (.A(_08093_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _14969_ (.A0(\rbzero.wall_tracer.stepDistX[-10] ),
    .A1(_07892_),
    .S(_08092_),
    .X(_08094_));
 sky130_fd_sc_hd__clkbuf_1 _14970_ (.A(_08094_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _14971_ (.A0(\rbzero.wall_tracer.stepDistX[-9] ),
    .A1(_07907_),
    .S(_08092_),
    .X(_08095_));
 sky130_fd_sc_hd__clkbuf_1 _14972_ (.A(_08095_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _14973_ (.A0(\rbzero.wall_tracer.stepDistX[-8] ),
    .A1(_07923_),
    .S(_08092_),
    .X(_08096_));
 sky130_fd_sc_hd__clkbuf_1 _14974_ (.A(_08096_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _14975_ (.A0(\rbzero.wall_tracer.stepDistX[-7] ),
    .A1(_07935_),
    .S(_08092_),
    .X(_08097_));
 sky130_fd_sc_hd__clkbuf_1 _14976_ (.A(_08097_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _14977_ (.A0(\rbzero.wall_tracer.stepDistX[-6] ),
    .A1(_07944_),
    .S(_08092_),
    .X(_08098_));
 sky130_fd_sc_hd__clkbuf_1 _14978_ (.A(_08098_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _14979_ (.A0(\rbzero.wall_tracer.stepDistX[-5] ),
    .A1(_07954_),
    .S(_08092_),
    .X(_08099_));
 sky130_fd_sc_hd__clkbuf_1 _14980_ (.A(_08099_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _14981_ (.A0(\rbzero.wall_tracer.stepDistX[-4] ),
    .A1(_07964_),
    .S(_08092_),
    .X(_08100_));
 sky130_fd_sc_hd__clkbuf_1 _14982_ (.A(_08100_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _14983_ (.A0(\rbzero.wall_tracer.stepDistX[-3] ),
    .A1(_07971_),
    .S(_08092_),
    .X(_08101_));
 sky130_fd_sc_hd__clkbuf_1 _14984_ (.A(_08101_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _14985_ (.A0(\rbzero.wall_tracer.stepDistX[-2] ),
    .A1(_07975_),
    .S(_08092_),
    .X(_08102_));
 sky130_fd_sc_hd__clkbuf_1 _14986_ (.A(_08102_),
    .X(_00444_));
 sky130_fd_sc_hd__buf_4 _14987_ (.A(_08091_),
    .X(_08103_));
 sky130_fd_sc_hd__mux2_1 _14988_ (.A0(\rbzero.wall_tracer.stepDistX[-1] ),
    .A1(_07982_),
    .S(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__clkbuf_1 _14989_ (.A(_08104_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _14990_ (.A0(\rbzero.wall_tracer.stepDistX[0] ),
    .A1(_07992_),
    .S(_08103_),
    .X(_08105_));
 sky130_fd_sc_hd__clkbuf_1 _14991_ (.A(_08105_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _14992_ (.A0(\rbzero.wall_tracer.stepDistX[1] ),
    .A1(_07996_),
    .S(_08103_),
    .X(_08106_));
 sky130_fd_sc_hd__clkbuf_1 _14993_ (.A(_08106_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _14994_ (.A0(\rbzero.wall_tracer.stepDistX[2] ),
    .A1(_08000_),
    .S(_08103_),
    .X(_08107_));
 sky130_fd_sc_hd__clkbuf_1 _14995_ (.A(_08107_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _14996_ (.A0(\rbzero.wall_tracer.stepDistX[3] ),
    .A1(_08006_),
    .S(_08103_),
    .X(_08108_));
 sky130_fd_sc_hd__clkbuf_1 _14997_ (.A(_08108_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _14998_ (.A0(\rbzero.wall_tracer.stepDistX[4] ),
    .A1(_08012_),
    .S(_08103_),
    .X(_08109_));
 sky130_fd_sc_hd__clkbuf_1 _14999_ (.A(_08109_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _15000_ (.A0(\rbzero.wall_tracer.stepDistX[5] ),
    .A1(_08015_),
    .S(_08103_),
    .X(_08110_));
 sky130_fd_sc_hd__clkbuf_1 _15001_ (.A(_08110_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _15002_ (.A0(\rbzero.wall_tracer.stepDistX[6] ),
    .A1(_08018_),
    .S(_08103_),
    .X(_08111_));
 sky130_fd_sc_hd__clkbuf_1 _15003_ (.A(_08111_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _15004_ (.A0(\rbzero.wall_tracer.stepDistX[7] ),
    .A1(_08023_),
    .S(_08103_),
    .X(_08112_));
 sky130_fd_sc_hd__clkbuf_1 _15005_ (.A(_08112_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _15006_ (.A0(\rbzero.wall_tracer.stepDistX[8] ),
    .A1(_08027_),
    .S(_08103_),
    .X(_08113_));
 sky130_fd_sc_hd__clkbuf_1 _15007_ (.A(_08113_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _15008_ (.A0(\rbzero.wall_tracer.stepDistX[9] ),
    .A1(_08029_),
    .S(_08091_),
    .X(_08114_));
 sky130_fd_sc_hd__clkbuf_1 _15009_ (.A(_08114_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _15010_ (.A0(\rbzero.wall_tracer.stepDistX[10] ),
    .A1(_08031_),
    .S(_08091_),
    .X(_08115_));
 sky130_fd_sc_hd__clkbuf_1 _15011_ (.A(_08115_),
    .X(_00456_));
 sky130_fd_sc_hd__buf_4 _15012_ (.A(_03974_),
    .X(_08116_));
 sky130_fd_sc_hd__clkbuf_4 _15013_ (.A(_08116_),
    .X(_08117_));
 sky130_fd_sc_hd__and2_1 _15014_ (.A(_08117_),
    .B(_05057_),
    .X(_08118_));
 sky130_fd_sc_hd__clkbuf_1 _15015_ (.A(_08118_),
    .X(_00457_));
 sky130_fd_sc_hd__nor2_1 _15016_ (.A(net63),
    .B(_05297_),
    .Y(_00458_));
 sky130_fd_sc_hd__and2_1 _15017_ (.A(_08117_),
    .B(_05382_),
    .X(_08119_));
 sky130_fd_sc_hd__clkbuf_1 _15018_ (.A(_08119_),
    .X(_00459_));
 sky130_fd_sc_hd__and2_1 _15019_ (.A(_08117_),
    .B(_05470_),
    .X(_08120_));
 sky130_fd_sc_hd__clkbuf_1 _15020_ (.A(_08120_),
    .X(_00460_));
 sky130_fd_sc_hd__and2_1 _15021_ (.A(_08117_),
    .B(_05551_),
    .X(_08121_));
 sky130_fd_sc_hd__clkbuf_1 _15022_ (.A(_08121_),
    .X(_00461_));
 sky130_fd_sc_hd__and2_1 _15023_ (.A(_08117_),
    .B(_05632_),
    .X(_08122_));
 sky130_fd_sc_hd__clkbuf_1 _15024_ (.A(_08122_),
    .X(_00462_));
 sky130_fd_sc_hd__buf_8 _15025_ (.A(_06106_),
    .X(_08123_));
 sky130_fd_sc_hd__buf_6 _15026_ (.A(_08123_),
    .X(_08124_));
 sky130_fd_sc_hd__nand2_1 _15027_ (.A(_08124_),
    .B(_08033_),
    .Y(_08125_));
 sky130_fd_sc_hd__nor2_1 _15028_ (.A(_06142_),
    .B(_06248_),
    .Y(_08126_));
 sky130_fd_sc_hd__or3_1 _15029_ (.A(_06159_),
    .B(_06233_),
    .C(_08126_),
    .X(_08127_));
 sky130_fd_sc_hd__a21bo_1 _15030_ (.A1(\rbzero.mapdyw[0] ),
    .A2(_06159_),
    .B1_N(_08127_),
    .X(_08128_));
 sky130_fd_sc_hd__mux2_1 _15031_ (.A0(_08128_),
    .A1(\rbzero.mapdxw[0] ),
    .S(_06151_),
    .X(_08129_));
 sky130_fd_sc_hd__a21o_1 _15032_ (.A1(_08124_),
    .A2(_08033_),
    .B1(\rbzero.wall_hot[0] ),
    .X(_08130_));
 sky130_fd_sc_hd__o211a_1 _15033_ (.A1(_08125_),
    .A2(_08129_),
    .B1(_08130_),
    .C1(_08085_),
    .X(_00463_));
 sky130_fd_sc_hd__nor2_1 _15034_ (.A(_06159_),
    .B(_08126_),
    .Y(_08131_));
 sky130_fd_sc_hd__a22o_1 _15035_ (.A1(\rbzero.mapdyw[1] ),
    .A2(_06159_),
    .B1(_06255_),
    .B2(_08131_),
    .X(_08132_));
 sky130_fd_sc_hd__mux2_1 _15036_ (.A0(_08132_),
    .A1(\rbzero.mapdxw[1] ),
    .S(_06151_),
    .X(_08133_));
 sky130_fd_sc_hd__buf_4 _15037_ (.A(_04432_),
    .X(_08134_));
 sky130_fd_sc_hd__buf_4 _15038_ (.A(_08134_),
    .X(_08135_));
 sky130_fd_sc_hd__buf_6 _15039_ (.A(_08135_),
    .X(_08136_));
 sky130_fd_sc_hd__a21oi_1 _15040_ (.A1(_04526_),
    .A2(_08125_),
    .B1(_08136_),
    .Y(_08137_));
 sky130_fd_sc_hd__o21a_1 _15041_ (.A1(_08125_),
    .A2(_08133_),
    .B1(_08137_),
    .X(_00464_));
 sky130_fd_sc_hd__buf_4 _15042_ (.A(_04464_),
    .X(_08138_));
 sky130_fd_sc_hd__nor2_1 _15043_ (.A(_06217_),
    .B(_08035_),
    .Y(_08139_));
 sky130_fd_sc_hd__a21oi_1 _15044_ (.A1(_08138_),
    .A2(_08035_),
    .B1(_08139_),
    .Y(_08140_));
 sky130_fd_sc_hd__nor2_1 _15045_ (.A(_08136_),
    .B(_08140_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _15046_ (.A(\rbzero.trace_state[3] ),
    .B(\rbzero.trace_state[2] ),
    .Y(_08141_));
 sky130_fd_sc_hd__nor2_1 _15047_ (.A(_04430_),
    .B(_08141_),
    .Y(_08142_));
 sky130_fd_sc_hd__clkbuf_4 _15048_ (.A(_08142_),
    .X(_08143_));
 sky130_fd_sc_hd__buf_4 _15049_ (.A(_08143_),
    .X(_08144_));
 sky130_fd_sc_hd__clkbuf_8 _15050_ (.A(_08144_),
    .X(_08145_));
 sky130_fd_sc_hd__or2_1 _15051_ (.A(_04430_),
    .B(_08141_),
    .X(_08146_));
 sky130_fd_sc_hd__clkbuf_4 _15052_ (.A(_08146_),
    .X(_08147_));
 sky130_fd_sc_hd__buf_4 _15053_ (.A(_08147_),
    .X(_08148_));
 sky130_fd_sc_hd__buf_6 _15054_ (.A(_06260_),
    .X(_08149_));
 sky130_fd_sc_hd__nand2_2 _15055_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08149_),
    .Y(_08150_));
 sky130_fd_sc_hd__clkbuf_4 _15056_ (.A(_08150_),
    .X(_08151_));
 sky130_fd_sc_hd__clkbuf_4 _15057_ (.A(_08151_),
    .X(_08152_));
 sky130_fd_sc_hd__mux2_1 _15058_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .S(_04463_),
    .X(_08153_));
 sky130_fd_sc_hd__or2_1 _15059_ (.A(_08147_),
    .B(_08153_),
    .X(_08154_));
 sky130_fd_sc_hd__and2_1 _15060_ (.A(\rbzero.trace_state[1] ),
    .B(_06259_),
    .X(_08155_));
 sky130_fd_sc_hd__nand2_4 _15061_ (.A(\rbzero.trace_state[0] ),
    .B(_08155_),
    .Y(_08156_));
 sky130_fd_sc_hd__buf_4 _15062_ (.A(_08156_),
    .X(_08157_));
 sky130_fd_sc_hd__buf_4 _15063_ (.A(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__o211a_2 _15064_ (.A1(_07892_),
    .A2(_08144_),
    .B1(_08154_),
    .C1(_08158_),
    .X(_08159_));
 sky130_fd_sc_hd__clkbuf_4 _15065_ (.A(_08155_),
    .X(_08160_));
 sky130_fd_sc_hd__clkbuf_8 _15066_ (.A(_08160_),
    .X(_08161_));
 sky130_fd_sc_hd__nor2_8 _15067_ (.A(\rbzero.trace_state[0] ),
    .B(_06260_),
    .Y(_08162_));
 sky130_fd_sc_hd__a21o_1 _15068_ (.A1(\rbzero.wall_tracer.stepDistY[-10] ),
    .A2(_08161_),
    .B1(_08162_),
    .X(_08163_));
 sky130_fd_sc_hd__nor2_2 _15069_ (.A(_08159_),
    .B(_08163_),
    .Y(_08164_));
 sky130_fd_sc_hd__nand2_4 _15070_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08149_),
    .Y(_08165_));
 sky130_fd_sc_hd__clkbuf_4 _15071_ (.A(_08165_),
    .X(_08166_));
 sky130_fd_sc_hd__mux2_1 _15072_ (.A0(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .S(_04463_),
    .X(_08167_));
 sky130_fd_sc_hd__and3_2 _15073_ (.A(_04436_),
    .B(\rbzero.trace_state[0] ),
    .C(_06259_),
    .X(_08168_));
 sky130_fd_sc_hd__a21o_1 _15074_ (.A1(_08144_),
    .A2(_08167_),
    .B1(_08168_),
    .X(_08169_));
 sky130_fd_sc_hd__a21o_1 _15075_ (.A1(_07867_),
    .A2(_08148_),
    .B1(_08169_),
    .X(_08170_));
 sky130_fd_sc_hd__o211ai_4 _15076_ (.A1(\rbzero.wall_tracer.stepDistY[-11] ),
    .A2(_08149_),
    .B1(_06262_),
    .C1(_08170_),
    .Y(_08171_));
 sky130_fd_sc_hd__or4_2 _15077_ (.A(_08152_),
    .B(_08164_),
    .C(_08166_),
    .D(_08171_),
    .X(_08172_));
 sky130_fd_sc_hd__o21ai_1 _15078_ (.A1(_07969_),
    .A2(_07970_),
    .B1(_08147_),
    .Y(_08173_));
 sky130_fd_sc_hd__nand2_1 _15079_ (.A(\rbzero.side_hot ),
    .B(_06353_),
    .Y(_08174_));
 sky130_fd_sc_hd__o211a_1 _15080_ (.A1(_04463_),
    .A2(_06053_),
    .B1(_08142_),
    .C1(_08174_),
    .X(_08175_));
 sky130_fd_sc_hd__nor2_1 _15081_ (.A(_08160_),
    .B(_08175_),
    .Y(_08176_));
 sky130_fd_sc_hd__a2bb2o_2 _15082_ (.A1_N(\rbzero.wall_tracer.stepDistY[-3] ),
    .A2_N(_08156_),
    .B1(_08173_),
    .B2(_08176_),
    .X(_08177_));
 sky130_fd_sc_hd__o21bai_4 _15083_ (.A1(\rbzero.wall_tracer.stepDistX[-3] ),
    .A2(_06262_),
    .B1_N(_08177_),
    .Y(_08178_));
 sky130_fd_sc_hd__nor4_1 _15084_ (.A(\rbzero.wall_tracer.rayAddendX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .C(_06375_),
    .D(_06366_),
    .Y(_08179_));
 sky130_fd_sc_hd__and4b_1 _15085_ (.A_N(_06389_),
    .B(_06362_),
    .C(_06382_),
    .D(_08179_),
    .X(_08180_));
 sky130_fd_sc_hd__and3_1 _15086_ (.A(_06353_),
    .B(_06358_),
    .C(_08180_),
    .X(_08181_));
 sky130_fd_sc_hd__and3_1 _15087_ (.A(_06402_),
    .B(_06349_),
    .C(_08181_),
    .X(_08182_));
 sky130_fd_sc_hd__nor2_1 _15088_ (.A(_06396_),
    .B(_06397_),
    .Y(_08183_));
 sky130_fd_sc_hd__nor2_1 _15089_ (.A(_06341_),
    .B(_08183_),
    .Y(_08184_));
 sky130_fd_sc_hd__a31o_2 _15090_ (.A1(_06335_),
    .A2(_08182_),
    .A3(_08184_),
    .B1(_06426_),
    .X(_08185_));
 sky130_fd_sc_hd__xnor2_1 _15091_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_08186_));
 sky130_fd_sc_hd__or2_1 _15092_ (.A(_08185_),
    .B(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__nand2_1 _15093_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(_08185_),
    .Y(_08188_));
 sky130_fd_sc_hd__xnor2_1 _15094_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .B(\rbzero.debug_overlay.playerY[-9] ),
    .Y(_08189_));
 sky130_fd_sc_hd__inv_2 _15095_ (.A(\rbzero.debug_overlay.playerY[-8] ),
    .Y(_08190_));
 sky130_fd_sc_hd__mux2_1 _15096_ (.A0(_08189_),
    .A1(_08190_),
    .S(_06075_),
    .X(_08191_));
 sky130_fd_sc_hd__nor2_1 _15097_ (.A(\rbzero.wall_tracer.visualWallDist[-8] ),
    .B(_08160_),
    .Y(_08192_));
 sky130_fd_sc_hd__mux2_1 _15098_ (.A0(_08191_),
    .A1(_08192_),
    .S(_08156_),
    .X(_08193_));
 sky130_fd_sc_hd__a31o_1 _15099_ (.A1(_08162_),
    .A2(_08187_),
    .A3(_08188_),
    .B1(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__buf_2 _15100_ (.A(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__a31o_1 _15101_ (.A1(_07866_),
    .A2(_07958_),
    .A3(_07963_),
    .B1(_08143_),
    .X(_08196_));
 sky130_fd_sc_hd__nand2_1 _15102_ (.A(\rbzero.side_hot ),
    .B(_06358_),
    .Y(_08197_));
 sky130_fd_sc_hd__o211a_1 _15103_ (.A1(_04463_),
    .A2(_06056_),
    .B1(_08143_),
    .C1(_08197_),
    .X(_08198_));
 sky130_fd_sc_hd__nor2_1 _15104_ (.A(_08160_),
    .B(_08198_),
    .Y(_08199_));
 sky130_fd_sc_hd__a2bb2o_1 _15105_ (.A1_N(\rbzero.wall_tracer.stepDistY[-4] ),
    .A2_N(_08157_),
    .B1(_08196_),
    .B2(_08199_),
    .X(_08200_));
 sky130_fd_sc_hd__o21bai_4 _15106_ (.A1(\rbzero.wall_tracer.stepDistX[-4] ),
    .A2(_06262_),
    .B1_N(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__or3_1 _15107_ (.A(\rbzero.debug_overlay.playerY[-7] ),
    .B(\rbzero.debug_overlay.playerY[-8] ),
    .C(\rbzero.debug_overlay.playerY[-9] ),
    .X(_08202_));
 sky130_fd_sc_hd__o21ai_1 _15108_ (.A1(\rbzero.debug_overlay.playerY[-8] ),
    .A2(\rbzero.debug_overlay.playerY[-9] ),
    .B1(\rbzero.debug_overlay.playerY[-7] ),
    .Y(_08203_));
 sky130_fd_sc_hd__and2_1 _15109_ (.A(_08202_),
    .B(_08203_),
    .X(_08204_));
 sky130_fd_sc_hd__mux2_1 _15110_ (.A0(_08204_),
    .A1(\rbzero.debug_overlay.playerY[-7] ),
    .S(_06075_),
    .X(_08205_));
 sky130_fd_sc_hd__mux2_1 _15111_ (.A0(\rbzero.wall_tracer.visualWallDist[-7] ),
    .A1(_08205_),
    .S(_08168_),
    .X(_08206_));
 sky130_fd_sc_hd__or3_1 _15112_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .B(\rbzero.debug_overlay.playerX[-8] ),
    .C(\rbzero.debug_overlay.playerX[-9] ),
    .X(_08207_));
 sky130_fd_sc_hd__o21ai_1 _15113_ (.A1(\rbzero.debug_overlay.playerX[-8] ),
    .A2(\rbzero.debug_overlay.playerX[-9] ),
    .B1(\rbzero.debug_overlay.playerX[-7] ),
    .Y(_08208_));
 sky130_fd_sc_hd__nand2_1 _15114_ (.A(_08207_),
    .B(_08208_),
    .Y(_08209_));
 sky130_fd_sc_hd__nor2_1 _15115_ (.A(_08185_),
    .B(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__a211o_1 _15116_ (.A1(\rbzero.debug_overlay.playerX[-7] ),
    .A2(_08185_),
    .B1(_08210_),
    .C1(_06261_),
    .X(_08211_));
 sky130_fd_sc_hd__o21ai_2 _15117_ (.A1(_08162_),
    .A2(_08206_),
    .B1(_08211_),
    .Y(_08212_));
 sky130_fd_sc_hd__buf_2 _15118_ (.A(_08212_),
    .X(_08213_));
 sky130_fd_sc_hd__o22ai_1 _15119_ (.A1(_08178_),
    .A2(_08195_),
    .B1(_08201_),
    .B2(_08213_),
    .Y(_08214_));
 sky130_fd_sc_hd__or2_1 _15120_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_08207_),
    .X(_08215_));
 sky130_fd_sc_hd__nand2_1 _15121_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .B(_08207_),
    .Y(_08216_));
 sky130_fd_sc_hd__and2_1 _15122_ (.A(_08215_),
    .B(_08216_),
    .X(_08217_));
 sky130_fd_sc_hd__buf_4 _15123_ (.A(_08185_),
    .X(_08218_));
 sky130_fd_sc_hd__mux2_1 _15124_ (.A0(_08217_),
    .A1(\rbzero.debug_overlay.playerX[-6] ),
    .S(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__inv_2 _15125_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .Y(_08220_));
 sky130_fd_sc_hd__or2_1 _15126_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_08202_),
    .X(_08221_));
 sky130_fd_sc_hd__nand2_1 _15127_ (.A(\rbzero.debug_overlay.playerY[-6] ),
    .B(_08202_),
    .Y(_08222_));
 sky130_fd_sc_hd__nand2_1 _15128_ (.A(_08221_),
    .B(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__a31o_1 _15129_ (.A1(_06034_),
    .A2(_06074_),
    .A3(_08223_),
    .B1(_08157_),
    .X(_08224_));
 sky130_fd_sc_hd__a21oi_1 _15130_ (.A1(_08220_),
    .A2(_06076_),
    .B1(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__a211o_1 _15131_ (.A1(\rbzero.wall_tracer.visualWallDist[-6] ),
    .A2(_08158_),
    .B1(_08225_),
    .C1(_08162_),
    .X(_08226_));
 sky130_fd_sc_hd__o21ai_4 _15132_ (.A1(_06262_),
    .A2(_08219_),
    .B1(_08226_),
    .Y(_08227_));
 sky130_fd_sc_hd__buf_2 _15133_ (.A(_08227_),
    .X(_08228_));
 sky130_fd_sc_hd__nor2_2 _15134_ (.A(\rbzero.wall_tracer.stepDistX[-5] ),
    .B(_06261_),
    .Y(_08229_));
 sky130_fd_sc_hd__nand2_1 _15135_ (.A(\rbzero.side_hot ),
    .B(_06362_),
    .Y(_08230_));
 sky130_fd_sc_hd__o211a_1 _15136_ (.A1(\rbzero.side_hot ),
    .A2(_06058_),
    .B1(_08142_),
    .C1(_08230_),
    .X(_08231_));
 sky130_fd_sc_hd__a211o_1 _15137_ (.A1(_07954_),
    .A2(_08147_),
    .B1(_08231_),
    .C1(_08160_),
    .X(_08232_));
 sky130_fd_sc_hd__o21ai_4 _15138_ (.A1(\rbzero.wall_tracer.stepDistY[-5] ),
    .A2(_08157_),
    .B1(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__or2_1 _15139_ (.A(_08229_),
    .B(_08233_),
    .X(_08234_));
 sky130_fd_sc_hd__clkbuf_4 _15140_ (.A(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__nor2_1 _15141_ (.A(_08228_),
    .B(_08235_),
    .Y(_08236_));
 sky130_fd_sc_hd__or4_1 _15142_ (.A(_08178_),
    .B(_08213_),
    .C(_08195_),
    .D(_08201_),
    .X(_08237_));
 sky130_fd_sc_hd__a21bo_1 _15143_ (.A1(_08214_),
    .A2(_08236_),
    .B1_N(_08237_),
    .X(_08238_));
 sky130_fd_sc_hd__xor2_1 _15144_ (.A(\rbzero.debug_overlay.playerX[-5] ),
    .B(_08215_),
    .X(_08239_));
 sky130_fd_sc_hd__mux2_1 _15145_ (.A0(_08239_),
    .A1(\rbzero.debug_overlay.playerX[-5] ),
    .S(_08218_),
    .X(_08240_));
 sky130_fd_sc_hd__xor2_1 _15146_ (.A(\rbzero.debug_overlay.playerY[-5] ),
    .B(_08221_),
    .X(_08241_));
 sky130_fd_sc_hd__mux2_1 _15147_ (.A0(_08241_),
    .A1(\rbzero.debug_overlay.playerY[-5] ),
    .S(_06076_),
    .X(_08242_));
 sky130_fd_sc_hd__or2_1 _15148_ (.A(\rbzero.wall_tracer.visualWallDist[-5] ),
    .B(_08160_),
    .X(_08243_));
 sky130_fd_sc_hd__mux2_1 _15149_ (.A0(_08242_),
    .A1(_08243_),
    .S(_08157_),
    .X(_08244_));
 sky130_fd_sc_hd__o21ai_4 _15150_ (.A1(_06262_),
    .A2(_08240_),
    .B1(_08244_),
    .Y(_08245_));
 sky130_fd_sc_hd__buf_2 _15151_ (.A(_08245_),
    .X(_08246_));
 sky130_fd_sc_hd__o31ai_2 _15152_ (.A1(_07891_),
    .A2(_07942_),
    .A3(_07943_),
    .B1(_08147_),
    .Y(_08247_));
 sky130_fd_sc_hd__mux2_1 _15153_ (.A0(_06062_),
    .A1(_06389_),
    .S(_04463_),
    .X(_08248_));
 sky130_fd_sc_hd__a21oi_1 _15154_ (.A1(_08143_),
    .A2(_08248_),
    .B1(_08160_),
    .Y(_08249_));
 sky130_fd_sc_hd__a2bb2o_2 _15155_ (.A1_N(\rbzero.wall_tracer.stepDistY[-6] ),
    .A2_N(_08157_),
    .B1(_08247_),
    .B2(_08249_),
    .X(_08250_));
 sky130_fd_sc_hd__or2_1 _15156_ (.A(\rbzero.wall_tracer.stepDistX[-6] ),
    .B(_06261_),
    .X(_08251_));
 sky130_fd_sc_hd__or2b_1 _15157_ (.A(_08250_),
    .B_N(_08251_),
    .X(_08252_));
 sky130_fd_sc_hd__buf_2 _15158_ (.A(_08252_),
    .X(_08253_));
 sky130_fd_sc_hd__or3_1 _15159_ (.A(\rbzero.debug_overlay.playerX[-4] ),
    .B(\rbzero.debug_overlay.playerX[-5] ),
    .C(_08215_),
    .X(_08254_));
 sky130_fd_sc_hd__o21ai_1 _15160_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_08215_),
    .B1(\rbzero.debug_overlay.playerX[-4] ),
    .Y(_08255_));
 sky130_fd_sc_hd__and2_1 _15161_ (.A(_08254_),
    .B(_08255_),
    .X(_08256_));
 sky130_fd_sc_hd__mux2_1 _15162_ (.A0(_08256_),
    .A1(\rbzero.debug_overlay.playerX[-4] ),
    .S(_08185_),
    .X(_08257_));
 sky130_fd_sc_hd__inv_2 _15163_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_08258_));
 sky130_fd_sc_hd__or3_1 _15164_ (.A(\rbzero.debug_overlay.playerY[-4] ),
    .B(\rbzero.debug_overlay.playerY[-5] ),
    .C(_08221_),
    .X(_08259_));
 sky130_fd_sc_hd__o21ai_1 _15165_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_08221_),
    .B1(\rbzero.debug_overlay.playerY[-4] ),
    .Y(_08260_));
 sky130_fd_sc_hd__nand2_1 _15166_ (.A(_08259_),
    .B(_08260_),
    .Y(_08261_));
 sky130_fd_sc_hd__a31o_1 _15167_ (.A1(_06034_),
    .A2(_06074_),
    .A3(_08261_),
    .B1(_08156_),
    .X(_08262_));
 sky130_fd_sc_hd__a21oi_1 _15168_ (.A1(_08258_),
    .A2(_06076_),
    .B1(_08262_),
    .Y(_08263_));
 sky130_fd_sc_hd__a211o_1 _15169_ (.A1(\rbzero.wall_tracer.visualWallDist[-4] ),
    .A2(_08157_),
    .B1(_08263_),
    .C1(_08162_),
    .X(_08264_));
 sky130_fd_sc_hd__o21ai_4 _15170_ (.A1(_06262_),
    .A2(_08257_),
    .B1(_08264_),
    .Y(_08265_));
 sky130_fd_sc_hd__or4_1 _15171_ (.A(_08235_),
    .B(_08246_),
    .C(_08253_),
    .D(_08265_),
    .X(_08266_));
 sky130_fd_sc_hd__o22ai_1 _15172_ (.A1(_08235_),
    .A2(_08246_),
    .B1(_08253_),
    .B2(_08265_),
    .Y(_08267_));
 sky130_fd_sc_hd__nand2_1 _15173_ (.A(_08266_),
    .B(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__nor2_1 _15174_ (.A(\rbzero.wall_tracer.stepDistX[-7] ),
    .B(_06262_),
    .Y(_08269_));
 sky130_fd_sc_hd__a21o_1 _15175_ (.A1(_07933_),
    .A2(_07934_),
    .B1(_08143_),
    .X(_08270_));
 sky130_fd_sc_hd__nand2_1 _15176_ (.A(_04463_),
    .B(_06382_),
    .Y(_08271_));
 sky130_fd_sc_hd__o211a_1 _15177_ (.A1(_04463_),
    .A2(_06063_),
    .B1(_08143_),
    .C1(_08271_),
    .X(_08272_));
 sky130_fd_sc_hd__nor2_1 _15178_ (.A(_08160_),
    .B(_08272_),
    .Y(_08273_));
 sky130_fd_sc_hd__a2bb2o_4 _15179_ (.A1_N(\rbzero.wall_tracer.stepDistY[-7] ),
    .A2_N(_08157_),
    .B1(_08270_),
    .B2(_08273_),
    .X(_08274_));
 sky130_fd_sc_hd__or2_1 _15180_ (.A(_08269_),
    .B(_08274_),
    .X(_08275_));
 sky130_fd_sc_hd__clkbuf_4 _15181_ (.A(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__or2_1 _15182_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_08254_),
    .X(_08277_));
 sky130_fd_sc_hd__nand2_1 _15183_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .B(_08254_),
    .Y(_08278_));
 sky130_fd_sc_hd__and2_1 _15184_ (.A(_08277_),
    .B(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__mux2_1 _15185_ (.A0(_08279_),
    .A1(\rbzero.debug_overlay.playerX[-3] ),
    .S(_08218_),
    .X(_08280_));
 sky130_fd_sc_hd__or2_1 _15186_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_08259_),
    .X(_08281_));
 sky130_fd_sc_hd__nand2_1 _15187_ (.A(\rbzero.debug_overlay.playerY[-3] ),
    .B(_08259_),
    .Y(_08282_));
 sky130_fd_sc_hd__and2_1 _15188_ (.A(_08281_),
    .B(_08282_),
    .X(_08283_));
 sky130_fd_sc_hd__mux2_1 _15189_ (.A0(_08283_),
    .A1(\rbzero.debug_overlay.playerY[-3] ),
    .S(_06076_),
    .X(_08284_));
 sky130_fd_sc_hd__or2_1 _15190_ (.A(\rbzero.wall_tracer.visualWallDist[-3] ),
    .B(_08161_),
    .X(_08285_));
 sky130_fd_sc_hd__mux2_1 _15191_ (.A0(_08284_),
    .A1(_08285_),
    .S(_08158_),
    .X(_08286_));
 sky130_fd_sc_hd__o21ai_4 _15192_ (.A1(_06263_),
    .A2(_08280_),
    .B1(_08286_),
    .Y(_08287_));
 sky130_fd_sc_hd__nor2_1 _15193_ (.A(_08276_),
    .B(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__xnor2_1 _15194_ (.A(_08268_),
    .B(_08288_),
    .Y(_08289_));
 sky130_fd_sc_hd__xnor2_1 _15195_ (.A(_08238_),
    .B(_08289_),
    .Y(_08290_));
 sky130_fd_sc_hd__o22ai_1 _15196_ (.A1(_08246_),
    .A2(_08253_),
    .B1(_08265_),
    .B2(_08276_),
    .Y(_08291_));
 sky130_fd_sc_hd__inv_2 _15197_ (.A(\rbzero.wall_tracer.stepDistX[-8] ),
    .Y(_08292_));
 sky130_fd_sc_hd__a21o_1 _15198_ (.A1(_07919_),
    .A2(_07922_),
    .B1(_08143_),
    .X(_08293_));
 sky130_fd_sc_hd__mux2_1 _15199_ (.A0(_06065_),
    .A1(_06366_),
    .S(\rbzero.side_hot ),
    .X(_08294_));
 sky130_fd_sc_hd__a21oi_1 _15200_ (.A1(_08143_),
    .A2(_08294_),
    .B1(_08160_),
    .Y(_08295_));
 sky130_fd_sc_hd__a2bb2o_4 _15201_ (.A1_N(\rbzero.wall_tracer.stepDistY[-8] ),
    .A2_N(_08157_),
    .B1(_08293_),
    .B2(_08295_),
    .X(_08296_));
 sky130_fd_sc_hd__a21o_1 _15202_ (.A1(_08292_),
    .A2(_08162_),
    .B1(_08296_),
    .X(_08297_));
 sky130_fd_sc_hd__clkbuf_4 _15203_ (.A(_08297_),
    .X(_08298_));
 sky130_fd_sc_hd__nor2_1 _15204_ (.A(_08287_),
    .B(_08298_),
    .Y(_08299_));
 sky130_fd_sc_hd__or4_1 _15205_ (.A(_08245_),
    .B(_08252_),
    .C(_08265_),
    .D(_08275_),
    .X(_08300_));
 sky130_fd_sc_hd__a21bo_1 _15206_ (.A1(_08291_),
    .A2(_08299_),
    .B1_N(_08300_),
    .X(_08301_));
 sky130_fd_sc_hd__or2b_1 _15207_ (.A(_08290_),
    .B_N(_08301_),
    .X(_08302_));
 sky130_fd_sc_hd__a21bo_1 _15208_ (.A1(_08238_),
    .A2(_08289_),
    .B1_N(_08302_),
    .X(_08303_));
 sky130_fd_sc_hd__clkbuf_4 _15209_ (.A(_08164_),
    .X(_08304_));
 sky130_fd_sc_hd__o22ai_2 _15210_ (.A1(_08152_),
    .A2(_08304_),
    .B1(_08166_),
    .B2(_08171_),
    .Y(_08305_));
 sky130_fd_sc_hd__nand2_1 _15211_ (.A(_08172_),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__xor2_1 _15212_ (.A(\rbzero.debug_overlay.playerX[-2] ),
    .B(_08277_),
    .X(_08307_));
 sky130_fd_sc_hd__mux2_1 _15213_ (.A0(_08307_),
    .A1(\rbzero.debug_overlay.playerX[-2] ),
    .S(_08218_),
    .X(_08308_));
 sky130_fd_sc_hd__xor2_1 _15214_ (.A(\rbzero.debug_overlay.playerY[-2] ),
    .B(_08281_),
    .X(_08309_));
 sky130_fd_sc_hd__mux2_1 _15215_ (.A0(_08309_),
    .A1(\rbzero.debug_overlay.playerY[-2] ),
    .S(_06076_),
    .X(_08310_));
 sky130_fd_sc_hd__or2_1 _15216_ (.A(\rbzero.wall_tracer.visualWallDist[-2] ),
    .B(_08160_),
    .X(_08311_));
 sky130_fd_sc_hd__mux2_1 _15217_ (.A0(_08310_),
    .A1(_08311_),
    .S(_08158_),
    .X(_08312_));
 sky130_fd_sc_hd__o21ai_4 _15218_ (.A1(_06262_),
    .A2(_08308_),
    .B1(_08312_),
    .Y(_08313_));
 sky130_fd_sc_hd__or2_1 _15219_ (.A(_08298_),
    .B(_08313_),
    .X(_08314_));
 sky130_fd_sc_hd__or3_4 _15220_ (.A(\rbzero.debug_overlay.playerX[-1] ),
    .B(\rbzero.debug_overlay.playerX[-2] ),
    .C(_08277_),
    .X(_08315_));
 sky130_fd_sc_hd__o21ai_1 _15221_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_08277_),
    .B1(\rbzero.debug_overlay.playerX[-1] ),
    .Y(_08316_));
 sky130_fd_sc_hd__nand2_1 _15222_ (.A(_08315_),
    .B(_08316_),
    .Y(_08317_));
 sky130_fd_sc_hd__mux2_1 _15223_ (.A0(_08317_),
    .A1(_04692_),
    .S(_08218_),
    .X(_08318_));
 sky130_fd_sc_hd__nor2_1 _15224_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .B(_06087_),
    .Y(_08319_));
 sky130_fd_sc_hd__or3_2 _15225_ (.A(\rbzero.debug_overlay.playerY[-1] ),
    .B(\rbzero.debug_overlay.playerY[-2] ),
    .C(_08281_),
    .X(_08320_));
 sky130_fd_sc_hd__o21ai_1 _15226_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_08281_),
    .B1(\rbzero.debug_overlay.playerY[-1] ),
    .Y(_08321_));
 sky130_fd_sc_hd__nand2_1 _15227_ (.A(_08320_),
    .B(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__a31o_1 _15228_ (.A1(_06034_),
    .A2(_06074_),
    .A3(_08322_),
    .B1(_08158_),
    .X(_08323_));
 sky130_fd_sc_hd__o2bb2a_1 _15229_ (.A1_N(\rbzero.wall_tracer.visualWallDist[-1] ),
    .A2_N(_08158_),
    .B1(_08319_),
    .B2(_08323_),
    .X(_08324_));
 sky130_fd_sc_hd__mux2_4 _15230_ (.A0(_08318_),
    .A1(_08324_),
    .S(_06263_),
    .X(_08325_));
 sky130_fd_sc_hd__or3_1 _15231_ (.A(_08276_),
    .B(_08314_),
    .C(_08325_),
    .X(_08326_));
 sky130_fd_sc_hd__clkbuf_4 _15232_ (.A(_08325_),
    .X(_08327_));
 sky130_fd_sc_hd__buf_2 _15233_ (.A(_08313_),
    .X(_08328_));
 sky130_fd_sc_hd__nor2_1 _15234_ (.A(_08276_),
    .B(_08328_),
    .Y(_08329_));
 sky130_fd_sc_hd__o21bai_1 _15235_ (.A1(_08298_),
    .A2(_08327_),
    .B1_N(_08329_),
    .Y(_08330_));
 sky130_fd_sc_hd__nand2_1 _15236_ (.A(_08326_),
    .B(_08330_),
    .Y(_08331_));
 sky130_fd_sc_hd__nor2_1 _15237_ (.A(\rbzero.wall_tracer.stepDistX[-9] ),
    .B(_06262_),
    .Y(_08332_));
 sky130_fd_sc_hd__mux2_1 _15238_ (.A0(_06066_),
    .A1(_06375_),
    .S(_04463_),
    .X(_08333_));
 sky130_fd_sc_hd__mux2_1 _15239_ (.A0(_07907_),
    .A1(_08333_),
    .S(_08143_),
    .X(_08334_));
 sky130_fd_sc_hd__o22ai_4 _15240_ (.A1(\rbzero.wall_tracer.stepDistY[-9] ),
    .A2(_08157_),
    .B1(_08334_),
    .B2(_08161_),
    .Y(_08335_));
 sky130_fd_sc_hd__or2_1 _15241_ (.A(_08332_),
    .B(_08335_),
    .X(_08336_));
 sky130_fd_sc_hd__clkbuf_4 _15242_ (.A(_08336_),
    .X(_08337_));
 sky130_fd_sc_hd__clkbuf_8 _15243_ (.A(_08161_),
    .X(_08338_));
 sky130_fd_sc_hd__o32a_1 _15244_ (.A1(_06076_),
    .A2(_08158_),
    .A3(_08320_),
    .B1(_08338_),
    .B2(_08069_),
    .X(_08339_));
 sky130_fd_sc_hd__o31a_4 _15245_ (.A1(_06263_),
    .A2(_08218_),
    .A3(_08315_),
    .B1(_08339_),
    .X(_08340_));
 sky130_fd_sc_hd__or2_1 _15246_ (.A(_08337_),
    .B(_08340_),
    .X(_08341_));
 sky130_fd_sc_hd__xnor2_1 _15247_ (.A(_08331_),
    .B(_08341_),
    .Y(_08342_));
 sky130_fd_sc_hd__o22ai_4 _15248_ (.A1(\rbzero.wall_tracer.stepDistX[-10] ),
    .A2(_06263_),
    .B1(_08159_),
    .B2(_08163_),
    .Y(_08343_));
 sky130_fd_sc_hd__clkbuf_4 _15249_ (.A(_08343_),
    .X(_08344_));
 sky130_fd_sc_hd__nor2_1 _15250_ (.A(_08340_),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__nor2_1 _15251_ (.A(_08325_),
    .B(_08337_),
    .Y(_08346_));
 sky130_fd_sc_hd__xnor2_1 _15252_ (.A(_08314_),
    .B(_08346_),
    .Y(_08347_));
 sky130_fd_sc_hd__nand2_1 _15253_ (.A(_08345_),
    .B(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__o31a_1 _15254_ (.A1(_08314_),
    .A2(_08327_),
    .A3(_08337_),
    .B1(_08348_),
    .X(_08349_));
 sky130_fd_sc_hd__nor2_1 _15255_ (.A(_08342_),
    .B(_08349_),
    .Y(_08350_));
 sky130_fd_sc_hd__and2_1 _15256_ (.A(_08342_),
    .B(_08349_),
    .X(_08351_));
 sky130_fd_sc_hd__nor2_1 _15257_ (.A(_08350_),
    .B(_08351_),
    .Y(_08352_));
 sky130_fd_sc_hd__xnor2_1 _15258_ (.A(_08306_),
    .B(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__xnor2_1 _15259_ (.A(_08303_),
    .B(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__xnor2_1 _15260_ (.A(_08345_),
    .B(_08347_),
    .Y(_08355_));
 sky130_fd_sc_hd__nor2_1 _15261_ (.A(_08328_),
    .B(_08343_),
    .Y(_08356_));
 sky130_fd_sc_hd__buf_4 _15262_ (.A(_08162_),
    .X(_08357_));
 sky130_fd_sc_hd__a21boi_2 _15263_ (.A1(\rbzero.wall_tracer.stepDistX[-11] ),
    .A2(_08357_),
    .B1_N(_08171_),
    .Y(_08358_));
 sky130_fd_sc_hd__or2_1 _15264_ (.A(_08340_),
    .B(_08358_),
    .X(_08359_));
 sky130_fd_sc_hd__o22a_1 _15265_ (.A1(_08328_),
    .A2(_08337_),
    .B1(_08343_),
    .B2(_08325_),
    .X(_08360_));
 sky130_fd_sc_hd__o2bb2a_1 _15266_ (.A1_N(_08346_),
    .A2_N(_08356_),
    .B1(_08359_),
    .B2(_08360_),
    .X(_08361_));
 sky130_fd_sc_hd__xnor2_1 _15267_ (.A(_08355_),
    .B(_08361_),
    .Y(_08362_));
 sky130_fd_sc_hd__or3_2 _15268_ (.A(_08152_),
    .B(_08171_),
    .C(_08362_),
    .X(_08363_));
 sky130_fd_sc_hd__o21ai_1 _15269_ (.A1(_08355_),
    .A2(_08361_),
    .B1(_08363_),
    .Y(_08364_));
 sky130_fd_sc_hd__or2b_1 _15270_ (.A(_08354_),
    .B_N(_08364_),
    .X(_08365_));
 sky130_fd_sc_hd__a21boi_1 _15271_ (.A1(_08303_),
    .A2(_08353_),
    .B1_N(_08365_),
    .Y(_08366_));
 sky130_fd_sc_hd__or2_1 _15272_ (.A(_08172_),
    .B(_08366_),
    .X(_08367_));
 sky130_fd_sc_hd__buf_2 _15273_ (.A(_08178_),
    .X(_08368_));
 sky130_fd_sc_hd__buf_4 _15274_ (.A(_08246_),
    .X(_08369_));
 sky130_fd_sc_hd__clkbuf_4 _15275_ (.A(_08201_),
    .X(_08370_));
 sky130_fd_sc_hd__or2_1 _15276_ (.A(_08370_),
    .B(_08265_),
    .X(_08371_));
 sky130_fd_sc_hd__o21ai_1 _15277_ (.A1(_08368_),
    .A2(_08369_),
    .B1(_08371_),
    .Y(_08372_));
 sky130_fd_sc_hd__clkbuf_4 _15278_ (.A(_08287_),
    .X(_08373_));
 sky130_fd_sc_hd__nor2_1 _15279_ (.A(_08235_),
    .B(_08373_),
    .Y(_08374_));
 sky130_fd_sc_hd__or3_1 _15280_ (.A(_08368_),
    .B(_08246_),
    .C(_08371_),
    .X(_08375_));
 sky130_fd_sc_hd__a21bo_1 _15281_ (.A1(_08372_),
    .A2(_08374_),
    .B1_N(_08375_),
    .X(_08376_));
 sky130_fd_sc_hd__nor2_1 _15282_ (.A(_08368_),
    .B(_08265_),
    .Y(_08377_));
 sky130_fd_sc_hd__mux2_1 _15283_ (.A0(_06073_),
    .A1(_06349_),
    .S(\rbzero.side_hot ),
    .X(_08378_));
 sky130_fd_sc_hd__a21o_1 _15284_ (.A1(_08142_),
    .A2(_08378_),
    .B1(_08155_),
    .X(_08379_));
 sky130_fd_sc_hd__a21oi_2 _15285_ (.A1(_07975_),
    .A2(_08147_),
    .B1(_08379_),
    .Y(_08380_));
 sky130_fd_sc_hd__a21oi_1 _15286_ (.A1(\rbzero.wall_tracer.stepDistY[-2] ),
    .A2(_08168_),
    .B1(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__clkbuf_4 _15287_ (.A(_08381_),
    .X(_08382_));
 sky130_fd_sc_hd__a21boi_2 _15288_ (.A1(\rbzero.wall_tracer.stepDistX[-2] ),
    .A2(_08162_),
    .B1_N(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__clkbuf_4 _15289_ (.A(_08383_),
    .X(_08384_));
 sky130_fd_sc_hd__nor2_1 _15290_ (.A(_08246_),
    .B(_08384_),
    .Y(_08385_));
 sky130_fd_sc_hd__xnor2_1 _15291_ (.A(_08377_),
    .B(_08385_),
    .Y(_08386_));
 sky130_fd_sc_hd__or3_1 _15292_ (.A(_08370_),
    .B(_08373_),
    .C(_08386_),
    .X(_08387_));
 sky130_fd_sc_hd__o21ai_1 _15293_ (.A1(_08370_),
    .A2(_08373_),
    .B1(_08386_),
    .Y(_08388_));
 sky130_fd_sc_hd__nand2_1 _15294_ (.A(_08387_),
    .B(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__clkbuf_4 _15295_ (.A(_08195_),
    .X(_08390_));
 sky130_fd_sc_hd__inv_2 _15296_ (.A(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_08391_));
 sky130_fd_sc_hd__inv_2 _15297_ (.A(\rbzero.wall_tracer.stepDistY[0] ),
    .Y(_08392_));
 sky130_fd_sc_hd__or3b_2 _15298_ (.A(_06516_),
    .B(_07975_),
    .C_N(_07981_),
    .X(_08393_));
 sky130_fd_sc_hd__xor2_1 _15299_ (.A(_07992_),
    .B(_08393_),
    .X(_08394_));
 sky130_fd_sc_hd__inv_2 _15300_ (.A(\rbzero.side_hot ),
    .Y(_08395_));
 sky130_fd_sc_hd__a31o_1 _15301_ (.A1(_08395_),
    .A2(_06044_),
    .A3(_06045_),
    .B1(_08147_),
    .X(_08396_));
 sky130_fd_sc_hd__a21o_1 _15302_ (.A1(_04464_),
    .A2(_08183_),
    .B1(_08396_),
    .X(_08397_));
 sky130_fd_sc_hd__o21ai_2 _15303_ (.A1(_08144_),
    .A2(_08394_),
    .B1(_08397_),
    .Y(_08398_));
 sky130_fd_sc_hd__mux2_4 _15304_ (.A0(_08392_),
    .A1(_08398_),
    .S(_08158_),
    .X(_08399_));
 sky130_fd_sc_hd__mux2_2 _15305_ (.A0(_08391_),
    .A1(_08399_),
    .S(_06263_),
    .X(_08400_));
 sky130_fd_sc_hd__xor2_1 _15306_ (.A(_07975_),
    .B(_07982_),
    .X(_08401_));
 sky130_fd_sc_hd__nor2_1 _15307_ (.A(\rbzero.side_hot ),
    .B(_06055_),
    .Y(_08402_));
 sky130_fd_sc_hd__a211o_1 _15308_ (.A1(_04463_),
    .A2(_06402_),
    .B1(_08147_),
    .C1(_08402_),
    .X(_08403_));
 sky130_fd_sc_hd__o21a_2 _15309_ (.A1(_08143_),
    .A2(_08401_),
    .B1(_08403_),
    .X(_08404_));
 sky130_fd_sc_hd__buf_4 _15310_ (.A(_08168_),
    .X(_08405_));
 sky130_fd_sc_hd__nand2_1 _15311_ (.A(\rbzero.wall_tracer.stepDistY[-1] ),
    .B(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__nand2_1 _15312_ (.A(\rbzero.wall_tracer.stepDistX[-1] ),
    .B(_08357_),
    .Y(_08407_));
 sky130_fd_sc_hd__o211a_2 _15313_ (.A1(_08161_),
    .A2(_08404_),
    .B1(_08406_),
    .C1(_08407_),
    .X(_08408_));
 sky130_fd_sc_hd__clkbuf_4 _15314_ (.A(_08408_),
    .X(_08409_));
 sky130_fd_sc_hd__clkbuf_4 _15315_ (.A(_08213_),
    .X(_08410_));
 sky130_fd_sc_hd__o22a_1 _15316_ (.A1(_08390_),
    .A2(_08400_),
    .B1(_08409_),
    .B2(_08410_),
    .X(_08411_));
 sky130_fd_sc_hd__or2_1 _15317_ (.A(_08228_),
    .B(_08384_),
    .X(_08412_));
 sky130_fd_sc_hd__nor2_1 _15318_ (.A(_08410_),
    .B(_08400_),
    .Y(_08413_));
 sky130_fd_sc_hd__nor2_1 _15319_ (.A(_08390_),
    .B(_08409_),
    .Y(_08414_));
 sky130_fd_sc_hd__a2bb2o_1 _15320_ (.A1_N(_08411_),
    .A2_N(_08412_),
    .B1(_08413_),
    .B2(_08414_),
    .X(_08415_));
 sky130_fd_sc_hd__or2b_1 _15321_ (.A(_08389_),
    .B_N(_08415_),
    .X(_08416_));
 sky130_fd_sc_hd__or2b_1 _15322_ (.A(_08415_),
    .B_N(_08389_),
    .X(_08417_));
 sky130_fd_sc_hd__nand2_1 _15323_ (.A(_08416_),
    .B(_08417_),
    .Y(_08418_));
 sky130_fd_sc_hd__xnor2_1 _15324_ (.A(_08376_),
    .B(_08418_),
    .Y(_08419_));
 sky130_fd_sc_hd__inv_2 _15325_ (.A(\rbzero.wall_tracer.stepDistX[1] ),
    .Y(_08420_));
 sky130_fd_sc_hd__clkbuf_4 _15326_ (.A(_08158_),
    .X(_08421_));
 sky130_fd_sc_hd__inv_2 _15327_ (.A(\rbzero.wall_tracer.stepDistY[1] ),
    .Y(_08422_));
 sky130_fd_sc_hd__mux2_1 _15328_ (.A0(_06041_),
    .A1(_06341_),
    .S(_04464_),
    .X(_08423_));
 sky130_fd_sc_hd__nand2_1 _15329_ (.A(_08144_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__a21o_1 _15330_ (.A1(_07992_),
    .A2(_08393_),
    .B1(_07996_),
    .X(_08425_));
 sky130_fd_sc_hd__nand3_1 _15331_ (.A(_07992_),
    .B(_07996_),
    .C(_08393_),
    .Y(_08426_));
 sky130_fd_sc_hd__a21o_1 _15332_ (.A1(_08425_),
    .A2(_08426_),
    .B1(_08144_),
    .X(_08427_));
 sky130_fd_sc_hd__a21o_2 _15333_ (.A1(_08424_),
    .A2(_08427_),
    .B1(_08161_),
    .X(_08428_));
 sky130_fd_sc_hd__o221a_2 _15334_ (.A1(_08420_),
    .A2(_06263_),
    .B1(_08421_),
    .B2(_08422_),
    .C1(_08428_),
    .X(_08429_));
 sky130_fd_sc_hd__or4_1 _15335_ (.A(_08410_),
    .B(_08390_),
    .C(_08400_),
    .D(_08429_),
    .X(_08430_));
 sky130_fd_sc_hd__clkbuf_4 _15336_ (.A(_08390_),
    .X(_08431_));
 sky130_fd_sc_hd__o21bai_1 _15337_ (.A1(_08431_),
    .A2(_08429_),
    .B1_N(_08413_),
    .Y(_08432_));
 sky130_fd_sc_hd__nand2_1 _15338_ (.A(_08430_),
    .B(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__clkbuf_4 _15339_ (.A(_08228_),
    .X(_08434_));
 sky130_fd_sc_hd__nor2_1 _15340_ (.A(_08434_),
    .B(_08409_),
    .Y(_08435_));
 sky130_fd_sc_hd__xnor2_1 _15341_ (.A(_08433_),
    .B(_08435_),
    .Y(_08436_));
 sky130_fd_sc_hd__clkinv_2 _15342_ (.A(\rbzero.debug_overlay.playerY[-9] ),
    .Y(_08437_));
 sky130_fd_sc_hd__nor2_1 _15343_ (.A(_08437_),
    .B(_08158_),
    .Y(_08438_));
 sky130_fd_sc_hd__a221oi_2 _15344_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_06260_),
    .B1(_08162_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__buf_2 _15345_ (.A(_08439_),
    .X(_08440_));
 sky130_fd_sc_hd__clkbuf_4 _15346_ (.A(_08440_),
    .X(_08441_));
 sky130_fd_sc_hd__xor2_1 _15347_ (.A(_08000_),
    .B(_08425_),
    .X(_08442_));
 sky130_fd_sc_hd__nor2_1 _15348_ (.A(_04464_),
    .B(_06037_),
    .Y(_08443_));
 sky130_fd_sc_hd__a211o_1 _15349_ (.A1(_04464_),
    .A2(_06335_),
    .B1(_08147_),
    .C1(_08443_),
    .X(_08444_));
 sky130_fd_sc_hd__o21ai_4 _15350_ (.A1(_08144_),
    .A2(_08442_),
    .B1(_08444_),
    .Y(_08445_));
 sky130_fd_sc_hd__a22o_1 _15351_ (.A1(\rbzero.wall_tracer.stepDistX[2] ),
    .A2(_08357_),
    .B1(_08405_),
    .B2(\rbzero.wall_tracer.stepDistY[2] ),
    .X(_08446_));
 sky130_fd_sc_hd__a21oi_2 _15352_ (.A1(_08149_),
    .A2(_08445_),
    .B1(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__nor2_1 _15353_ (.A(_08441_),
    .B(_08447_),
    .Y(_08448_));
 sky130_fd_sc_hd__a2111o_1 _15354_ (.A1(_07992_),
    .A2(_08393_),
    .B1(_08006_),
    .C1(_08000_),
    .D1(_07996_),
    .X(_08449_));
 sky130_fd_sc_hd__buf_2 _15355_ (.A(_08449_),
    .X(_08450_));
 sky130_fd_sc_hd__o21ai_1 _15356_ (.A1(_08000_),
    .A2(_08425_),
    .B1(_08006_),
    .Y(_08451_));
 sky130_fd_sc_hd__nand2_1 _15357_ (.A(_04464_),
    .B(_06426_),
    .Y(_08452_));
 sky130_fd_sc_hd__or2_2 _15358_ (.A(_04464_),
    .B(_06034_),
    .X(_08453_));
 sky130_fd_sc_hd__a31o_2 _15359_ (.A1(_08144_),
    .A2(_08452_),
    .A3(_08453_),
    .B1(_08168_),
    .X(_08454_));
 sky130_fd_sc_hd__a31o_2 _15360_ (.A1(_08148_),
    .A2(_08450_),
    .A3(_08451_),
    .B1(_08454_),
    .X(_08455_));
 sky130_fd_sc_hd__nand2_1 _15361_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_06260_),
    .Y(_08456_));
 sky130_fd_sc_hd__buf_2 _15362_ (.A(_08456_),
    .X(_08457_));
 sky130_fd_sc_hd__buf_4 _15363_ (.A(_08457_),
    .X(_08458_));
 sky130_fd_sc_hd__nor2_2 _15364_ (.A(_08455_),
    .B(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__nand2_1 _15365_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08156_),
    .Y(_08460_));
 sky130_fd_sc_hd__buf_2 _15366_ (.A(_08460_),
    .X(_08461_));
 sky130_fd_sc_hd__nand2_1 _15367_ (.A(\rbzero.wall_tracer.stepDistY[4] ),
    .B(_08405_),
    .Y(_08462_));
 sky130_fd_sc_hd__nand2_1 _15368_ (.A(_08012_),
    .B(_08450_),
    .Y(_08463_));
 sky130_fd_sc_hd__or2_1 _15369_ (.A(_08011_),
    .B(_08450_),
    .X(_08464_));
 sky130_fd_sc_hd__a31o_1 _15370_ (.A1(_08148_),
    .A2(_08463_),
    .A3(_08464_),
    .B1(_08454_),
    .X(_08465_));
 sky130_fd_sc_hd__a21o_2 _15371_ (.A1(_08462_),
    .A2(_08465_),
    .B1(_08357_),
    .X(_08466_));
 sky130_fd_sc_hd__or2_1 _15372_ (.A(_08461_),
    .B(_08466_),
    .X(_08467_));
 sky130_fd_sc_hd__xnor2_1 _15373_ (.A(_08459_),
    .B(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__xnor2_2 _15374_ (.A(_08448_),
    .B(_08468_),
    .Y(_08469_));
 sky130_fd_sc_hd__or2_2 _15375_ (.A(_08429_),
    .B(_08440_),
    .X(_08470_));
 sky130_fd_sc_hd__nor2_2 _15376_ (.A(_08042_),
    .B(_08161_),
    .Y(_08471_));
 sky130_fd_sc_hd__nand2_1 _15377_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_06260_),
    .Y(_08472_));
 sky130_fd_sc_hd__buf_2 _15378_ (.A(_08472_),
    .X(_08473_));
 sky130_fd_sc_hd__o2bb2a_1 _15379_ (.A1_N(_08445_),
    .A2_N(_08471_),
    .B1(_08473_),
    .B2(_08455_),
    .X(_08474_));
 sky130_fd_sc_hd__buf_4 _15380_ (.A(_08149_),
    .X(_08475_));
 sky130_fd_sc_hd__nand2_1 _15381_ (.A(_08475_),
    .B(_08445_),
    .Y(_08476_));
 sky130_fd_sc_hd__or3b_1 _15382_ (.A(_08476_),
    .B(_08461_),
    .C_N(_08459_),
    .X(_08477_));
 sky130_fd_sc_hd__o21a_1 _15383_ (.A1(_08470_),
    .A2(_08474_),
    .B1(_08477_),
    .X(_08478_));
 sky130_fd_sc_hd__xor2_2 _15384_ (.A(_08469_),
    .B(_08478_),
    .X(_08479_));
 sky130_fd_sc_hd__xnor2_2 _15385_ (.A(_08436_),
    .B(_08479_),
    .Y(_08480_));
 sky130_fd_sc_hd__a21o_1 _15386_ (.A1(_08413_),
    .A2(_08414_),
    .B1(_08411_),
    .X(_08481_));
 sky130_fd_sc_hd__nor2_1 _15387_ (.A(_08434_),
    .B(_08384_),
    .Y(_08482_));
 sky130_fd_sc_hd__xnor2_1 _15388_ (.A(_08481_),
    .B(_08482_),
    .Y(_08483_));
 sky130_fd_sc_hd__nor2_2 _15389_ (.A(_08039_),
    .B(_08161_),
    .Y(_08484_));
 sky130_fd_sc_hd__a31oi_4 _15390_ (.A1(_08445_),
    .A2(_08484_),
    .A3(_08459_),
    .B1(_08474_),
    .Y(_08485_));
 sky130_fd_sc_hd__xor2_4 _15391_ (.A(_08470_),
    .B(_08485_),
    .X(_08486_));
 sky130_fd_sc_hd__or4b_1 _15392_ (.A(_08042_),
    .B(_08428_),
    .C(_08473_),
    .D_N(_08445_),
    .X(_08487_));
 sky130_fd_sc_hd__a2bb2o_1 _15393_ (.A1_N(_08042_),
    .A2_N(_08428_),
    .B1(_08445_),
    .B2(_08484_),
    .X(_08488_));
 sky130_fd_sc_hd__or4bb_1 _15394_ (.A(_08400_),
    .B(_08440_),
    .C_N(_08487_),
    .D_N(_08488_),
    .X(_08489_));
 sky130_fd_sc_hd__and2_1 _15395_ (.A(_08487_),
    .B(_08489_),
    .X(_08490_));
 sky130_fd_sc_hd__xor2_2 _15396_ (.A(_08486_),
    .B(_08490_),
    .X(_08491_));
 sky130_fd_sc_hd__nor2_1 _15397_ (.A(_08486_),
    .B(_08490_),
    .Y(_08492_));
 sky130_fd_sc_hd__a21o_1 _15398_ (.A1(_08483_),
    .A2(_08491_),
    .B1(_08492_),
    .X(_08493_));
 sky130_fd_sc_hd__xnor2_1 _15399_ (.A(_08480_),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__xnor2_1 _15400_ (.A(_08419_),
    .B(_08494_),
    .Y(_08495_));
 sky130_fd_sc_hd__xnor2_2 _15401_ (.A(_08483_),
    .B(_08491_),
    .Y(_08496_));
 sky130_fd_sc_hd__clkbuf_4 _15402_ (.A(_08400_),
    .X(_08497_));
 sky130_fd_sc_hd__a2bb2o_1 _15403_ (.A1_N(_08497_),
    .A2_N(_08441_),
    .B1(_08487_),
    .B2(_08488_),
    .X(_08498_));
 sky130_fd_sc_hd__and2_2 _15404_ (.A(_08424_),
    .B(_08427_),
    .X(_08499_));
 sky130_fd_sc_hd__o22ai_2 _15405_ (.A1(_08499_),
    .A2(_08473_),
    .B1(_08458_),
    .B2(_08399_),
    .Y(_08500_));
 sky130_fd_sc_hd__nor2_1 _15406_ (.A(_08408_),
    .B(_08440_),
    .Y(_08501_));
 sky130_fd_sc_hd__or3_2 _15407_ (.A(_08039_),
    .B(_08161_),
    .C(_08398_),
    .X(_08502_));
 sky130_fd_sc_hd__or3_1 _15408_ (.A(_08042_),
    .B(_08428_),
    .C(_08502_),
    .X(_08503_));
 sky130_fd_sc_hd__a21bo_1 _15409_ (.A1(_08500_),
    .A2(_08501_),
    .B1_N(_08503_),
    .X(_08504_));
 sky130_fd_sc_hd__nand3_1 _15410_ (.A(_08489_),
    .B(_08498_),
    .C(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__a21o_1 _15411_ (.A1(_08489_),
    .A2(_08498_),
    .B1(_08504_),
    .X(_08506_));
 sky130_fd_sc_hd__nor2_1 _15412_ (.A(_08195_),
    .B(_08384_),
    .Y(_08507_));
 sky130_fd_sc_hd__or3b_1 _15413_ (.A(_08410_),
    .B(_08408_),
    .C_N(_08507_),
    .X(_08508_));
 sky130_fd_sc_hd__o22ai_1 _15414_ (.A1(_08390_),
    .A2(_08409_),
    .B1(_08384_),
    .B2(_08410_),
    .Y(_08509_));
 sky130_fd_sc_hd__nand2_1 _15415_ (.A(_08508_),
    .B(_08509_),
    .Y(_08510_));
 sky130_fd_sc_hd__nor2_1 _15416_ (.A(_08368_),
    .B(_08228_),
    .Y(_08511_));
 sky130_fd_sc_hd__xnor2_1 _15417_ (.A(_08510_),
    .B(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__nand3_1 _15418_ (.A(_08505_),
    .B(_08506_),
    .C(_08512_),
    .Y(_08513_));
 sky130_fd_sc_hd__and2_1 _15419_ (.A(_08505_),
    .B(_08513_),
    .X(_08514_));
 sky130_fd_sc_hd__xor2_1 _15420_ (.A(_08496_),
    .B(_08514_),
    .X(_08515_));
 sky130_fd_sc_hd__clkbuf_4 _15421_ (.A(_08265_),
    .X(_08516_));
 sky130_fd_sc_hd__o22ai_1 _15422_ (.A1(_08370_),
    .A2(_08369_),
    .B1(_08516_),
    .B2(_08235_),
    .Y(_08517_));
 sky130_fd_sc_hd__nor2_1 _15423_ (.A(_08253_),
    .B(_08373_),
    .Y(_08518_));
 sky130_fd_sc_hd__or3_1 _15424_ (.A(_08235_),
    .B(_08246_),
    .C(_08371_),
    .X(_08519_));
 sky130_fd_sc_hd__a21bo_1 _15425_ (.A1(_08517_),
    .A2(_08518_),
    .B1_N(_08519_),
    .X(_08520_));
 sky130_fd_sc_hd__a21bo_1 _15426_ (.A1(_08509_),
    .A2(_08511_),
    .B1_N(_08508_),
    .X(_08521_));
 sky130_fd_sc_hd__and2_1 _15427_ (.A(_08375_),
    .B(_08372_),
    .X(_08522_));
 sky130_fd_sc_hd__xnor2_1 _15428_ (.A(_08522_),
    .B(_08374_),
    .Y(_08523_));
 sky130_fd_sc_hd__xor2_1 _15429_ (.A(_08521_),
    .B(_08523_),
    .X(_08524_));
 sky130_fd_sc_hd__xnor2_1 _15430_ (.A(_08520_),
    .B(_08524_),
    .Y(_08525_));
 sky130_fd_sc_hd__nor2_1 _15431_ (.A(_08496_),
    .B(_08514_),
    .Y(_08526_));
 sky130_fd_sc_hd__a21o_1 _15432_ (.A1(_08515_),
    .A2(_08525_),
    .B1(_08526_),
    .X(_08527_));
 sky130_fd_sc_hd__xnor2_1 _15433_ (.A(_08495_),
    .B(_08527_),
    .Y(_08528_));
 sky130_fd_sc_hd__and2b_1 _15434_ (.A_N(_08250_),
    .B(_08251_),
    .X(_08529_));
 sky130_fd_sc_hd__clkinv_2 _15435_ (.A(_08325_),
    .Y(_08530_));
 sky130_fd_sc_hd__o22a_1 _15436_ (.A1(_08253_),
    .A2(_08328_),
    .B1(_08325_),
    .B2(_08276_),
    .X(_08531_));
 sky130_fd_sc_hd__a31o_1 _15437_ (.A1(_08529_),
    .A2(_08530_),
    .A3(_08329_),
    .B1(_08531_),
    .X(_08532_));
 sky130_fd_sc_hd__or2_1 _15438_ (.A(_08298_),
    .B(_08340_),
    .X(_08533_));
 sky130_fd_sc_hd__xnor2_1 _15439_ (.A(_08532_),
    .B(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__clkbuf_4 _15440_ (.A(_08340_),
    .X(_08535_));
 sky130_fd_sc_hd__o31a_1 _15441_ (.A1(_08331_),
    .A2(_08337_),
    .A3(_08535_),
    .B1(_08326_),
    .X(_08536_));
 sky130_fd_sc_hd__nor2_1 _15442_ (.A(_08150_),
    .B(_08335_),
    .Y(_08537_));
 sky130_fd_sc_hd__o21ba_1 _15443_ (.A1(_08164_),
    .A2(_08165_),
    .B1_N(_08537_),
    .X(_08538_));
 sky130_fd_sc_hd__or3b_1 _15444_ (.A(_08164_),
    .B(_08165_),
    .C_N(_08537_),
    .X(_08539_));
 sky130_fd_sc_hd__and2b_1 _15445_ (.A_N(_08538_),
    .B(_08539_),
    .X(_08540_));
 sky130_fd_sc_hd__nand2_2 _15446_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08475_),
    .Y(_08541_));
 sky130_fd_sc_hd__or2_1 _15447_ (.A(_08171_),
    .B(_08541_),
    .X(_08542_));
 sky130_fd_sc_hd__xnor2_1 _15448_ (.A(_08540_),
    .B(_08542_),
    .Y(_08543_));
 sky130_fd_sc_hd__xor2_1 _15449_ (.A(_08534_),
    .B(_08536_),
    .X(_08544_));
 sky130_fd_sc_hd__nand2_1 _15450_ (.A(_08543_),
    .B(_08544_),
    .Y(_08545_));
 sky130_fd_sc_hd__o21ai_1 _15451_ (.A1(_08534_),
    .A2(_08536_),
    .B1(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__or2b_1 _15452_ (.A(_08523_),
    .B_N(_08521_),
    .X(_08547_));
 sky130_fd_sc_hd__or2b_1 _15453_ (.A(_08524_),
    .B_N(_08520_),
    .X(_08548_));
 sky130_fd_sc_hd__nor2_1 _15454_ (.A(_08165_),
    .B(_08335_),
    .Y(_08549_));
 sky130_fd_sc_hd__nor2_1 _15455_ (.A(_08151_),
    .B(_08296_),
    .Y(_08550_));
 sky130_fd_sc_hd__xnor2_1 _15456_ (.A(_08549_),
    .B(_08550_),
    .Y(_08551_));
 sky130_fd_sc_hd__or3_1 _15457_ (.A(_08304_),
    .B(_08541_),
    .C(_08551_),
    .X(_08552_));
 sky130_fd_sc_hd__clkbuf_4 _15458_ (.A(_08541_),
    .X(_08553_));
 sky130_fd_sc_hd__o21ai_1 _15459_ (.A1(_08304_),
    .A2(_08553_),
    .B1(_08551_),
    .Y(_08554_));
 sky130_fd_sc_hd__and2_1 _15460_ (.A(_08552_),
    .B(_08554_),
    .X(_08555_));
 sky130_fd_sc_hd__nor2_1 _15461_ (.A(_08253_),
    .B(_08328_),
    .Y(_08556_));
 sky130_fd_sc_hd__nor2_1 _15462_ (.A(_08235_),
    .B(_08327_),
    .Y(_08557_));
 sky130_fd_sc_hd__o22a_1 _15463_ (.A1(_08235_),
    .A2(_08328_),
    .B1(_08325_),
    .B2(_08253_),
    .X(_08558_));
 sky130_fd_sc_hd__a21o_1 _15464_ (.A1(_08556_),
    .A2(_08557_),
    .B1(_08558_),
    .X(_08559_));
 sky130_fd_sc_hd__or2_1 _15465_ (.A(_08276_),
    .B(_08340_),
    .X(_08560_));
 sky130_fd_sc_hd__xnor2_1 _15466_ (.A(_08559_),
    .B(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__or4_1 _15467_ (.A(_08253_),
    .B(_08276_),
    .C(_08328_),
    .D(_08327_),
    .X(_08562_));
 sky130_fd_sc_hd__o31a_1 _15468_ (.A1(_08298_),
    .A2(_08535_),
    .A3(_08531_),
    .B1(_08562_),
    .X(_08563_));
 sky130_fd_sc_hd__nor2_1 _15469_ (.A(_08561_),
    .B(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__and2_1 _15470_ (.A(_08561_),
    .B(_08563_),
    .X(_08565_));
 sky130_fd_sc_hd__nor2_1 _15471_ (.A(_08564_),
    .B(_08565_),
    .Y(_08566_));
 sky130_fd_sc_hd__xnor2_1 _15472_ (.A(_08555_),
    .B(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__a21o_1 _15473_ (.A1(_08547_),
    .A2(_08548_),
    .B1(_08567_),
    .X(_08568_));
 sky130_fd_sc_hd__nand3_1 _15474_ (.A(_08547_),
    .B(_08548_),
    .C(_08567_),
    .Y(_08569_));
 sky130_fd_sc_hd__nand2_1 _15475_ (.A(_08568_),
    .B(_08569_),
    .Y(_08570_));
 sky130_fd_sc_hd__xnor2_1 _15476_ (.A(_08546_),
    .B(_08570_),
    .Y(_08571_));
 sky130_fd_sc_hd__xnor2_1 _15477_ (.A(_08528_),
    .B(_08571_),
    .Y(_08572_));
 sky130_fd_sc_hd__xnor2_1 _15478_ (.A(_08515_),
    .B(_08525_),
    .Y(_08573_));
 sky130_fd_sc_hd__a21o_1 _15479_ (.A1(_08505_),
    .A2(_08506_),
    .B1(_08512_),
    .X(_08574_));
 sky130_fd_sc_hd__nand3_1 _15480_ (.A(_08503_),
    .B(_08500_),
    .C(_08501_),
    .Y(_08575_));
 sky130_fd_sc_hd__a21o_1 _15481_ (.A1(_08503_),
    .A2(_08500_),
    .B1(_08501_),
    .X(_08576_));
 sky130_fd_sc_hd__nor2_1 _15482_ (.A(_08404_),
    .B(_08457_),
    .Y(_08577_));
 sky130_fd_sc_hd__xnor2_2 _15483_ (.A(_08502_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__nor2_1 _15484_ (.A(_08383_),
    .B(_08440_),
    .Y(_08579_));
 sky130_fd_sc_hd__o21a_2 _15485_ (.A1(_08161_),
    .A2(_08404_),
    .B1(_08406_),
    .X(_08580_));
 sky130_fd_sc_hd__nand2_4 _15486_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_08156_),
    .Y(_08581_));
 sky130_fd_sc_hd__or3_1 _15487_ (.A(_08580_),
    .B(_08581_),
    .C(_08502_),
    .X(_08582_));
 sky130_fd_sc_hd__a21bo_1 _15488_ (.A1(_08578_),
    .A2(_08579_),
    .B1_N(_08582_),
    .X(_08583_));
 sky130_fd_sc_hd__a21o_1 _15489_ (.A1(_08575_),
    .A2(_08576_),
    .B1(_08583_),
    .X(_08584_));
 sky130_fd_sc_hd__nor2_1 _15490_ (.A(_08178_),
    .B(_08213_),
    .Y(_08585_));
 sky130_fd_sc_hd__xnor2_1 _15491_ (.A(_08585_),
    .B(_08507_),
    .Y(_08586_));
 sky130_fd_sc_hd__or3_1 _15492_ (.A(_08370_),
    .B(_08228_),
    .C(_08586_),
    .X(_08587_));
 sky130_fd_sc_hd__o21ai_1 _15493_ (.A1(_08370_),
    .A2(_08228_),
    .B1(_08586_),
    .Y(_08588_));
 sky130_fd_sc_hd__and2_1 _15494_ (.A(_08587_),
    .B(_08588_),
    .X(_08589_));
 sky130_fd_sc_hd__and3_1 _15495_ (.A(_08575_),
    .B(_08576_),
    .C(_08583_),
    .X(_08590_));
 sky130_fd_sc_hd__a21o_1 _15496_ (.A1(_08584_),
    .A2(_08589_),
    .B1(_08590_),
    .X(_08591_));
 sky130_fd_sc_hd__a21o_1 _15497_ (.A1(_08513_),
    .A2(_08574_),
    .B1(_08591_),
    .X(_08592_));
 sky130_fd_sc_hd__a21bo_1 _15498_ (.A1(_08267_),
    .A2(_08288_),
    .B1_N(_08266_),
    .X(_08593_));
 sky130_fd_sc_hd__a21bo_1 _15499_ (.A1(_08585_),
    .A2(_08507_),
    .B1_N(_08587_),
    .X(_08594_));
 sky130_fd_sc_hd__nand2_1 _15500_ (.A(_08519_),
    .B(_08517_),
    .Y(_08595_));
 sky130_fd_sc_hd__xor2_1 _15501_ (.A(_08595_),
    .B(_08518_),
    .X(_08596_));
 sky130_fd_sc_hd__xor2_1 _15502_ (.A(_08594_),
    .B(_08596_),
    .X(_08597_));
 sky130_fd_sc_hd__xnor2_1 _15503_ (.A(_08593_),
    .B(_08597_),
    .Y(_08598_));
 sky130_fd_sc_hd__nand3_1 _15504_ (.A(_08513_),
    .B(_08574_),
    .C(_08591_),
    .Y(_08599_));
 sky130_fd_sc_hd__a21boi_1 _15505_ (.A1(_08592_),
    .A2(_08598_),
    .B1_N(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__nor2_1 _15506_ (.A(_08573_),
    .B(_08600_),
    .Y(_08601_));
 sky130_fd_sc_hd__and2_1 _15507_ (.A(_08573_),
    .B(_08600_),
    .X(_08602_));
 sky130_fd_sc_hd__nor2_1 _15508_ (.A(_08601_),
    .B(_08602_),
    .Y(_08603_));
 sky130_fd_sc_hd__a31o_1 _15509_ (.A1(_08172_),
    .A2(_08305_),
    .A3(_08352_),
    .B1(_08350_),
    .X(_08604_));
 sky130_fd_sc_hd__or2b_1 _15510_ (.A(_08596_),
    .B_N(_08594_),
    .X(_08605_));
 sky130_fd_sc_hd__or2b_1 _15511_ (.A(_08597_),
    .B_N(_08593_),
    .X(_08606_));
 sky130_fd_sc_hd__or2_1 _15512_ (.A(_08543_),
    .B(_08544_),
    .X(_08607_));
 sky130_fd_sc_hd__nand2_1 _15513_ (.A(_08545_),
    .B(_08607_),
    .Y(_08608_));
 sky130_fd_sc_hd__a21o_1 _15514_ (.A1(_08605_),
    .A2(_08606_),
    .B1(_08608_),
    .X(_08609_));
 sky130_fd_sc_hd__nand3_1 _15515_ (.A(_08605_),
    .B(_08606_),
    .C(_08608_),
    .Y(_08610_));
 sky130_fd_sc_hd__nand2_1 _15516_ (.A(_08609_),
    .B(_08610_),
    .Y(_08611_));
 sky130_fd_sc_hd__xnor2_1 _15517_ (.A(_08604_),
    .B(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__a21oi_1 _15518_ (.A1(_08603_),
    .A2(_08612_),
    .B1(_08601_),
    .Y(_08613_));
 sky130_fd_sc_hd__xor2_1 _15519_ (.A(_08572_),
    .B(_08613_),
    .X(_08614_));
 sky130_fd_sc_hd__or2b_1 _15520_ (.A(_08611_),
    .B_N(_08604_),
    .X(_08615_));
 sky130_fd_sc_hd__buf_4 _15521_ (.A(_08171_),
    .X(_08616_));
 sky130_fd_sc_hd__nand2_4 _15522_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08149_),
    .Y(_08617_));
 sky130_fd_sc_hd__clkbuf_4 _15523_ (.A(_08617_),
    .X(_08618_));
 sky130_fd_sc_hd__or2_1 _15524_ (.A(_08616_),
    .B(_08618_),
    .X(_08619_));
 sky130_fd_sc_hd__clkbuf_4 _15525_ (.A(_08553_),
    .X(_08620_));
 sky130_fd_sc_hd__o31a_1 _15526_ (.A1(_08616_),
    .A2(_08538_),
    .A3(_08620_),
    .B1(_08539_),
    .X(_08621_));
 sky130_fd_sc_hd__nor2_1 _15527_ (.A(_08619_),
    .B(_08621_),
    .Y(_08622_));
 sky130_fd_sc_hd__and2_1 _15528_ (.A(_08619_),
    .B(_08621_),
    .X(_08623_));
 sky130_fd_sc_hd__or2_1 _15529_ (.A(_08622_),
    .B(_08623_),
    .X(_08624_));
 sky130_fd_sc_hd__a21oi_2 _15530_ (.A1(_08609_),
    .A2(_08615_),
    .B1(_08624_),
    .Y(_08625_));
 sky130_fd_sc_hd__and3_1 _15531_ (.A(_08609_),
    .B(_08615_),
    .C(_08624_),
    .X(_08626_));
 sky130_fd_sc_hd__nor2_1 _15532_ (.A(_08625_),
    .B(_08626_),
    .Y(_08627_));
 sky130_fd_sc_hd__xnor2_1 _15533_ (.A(_08614_),
    .B(_08627_),
    .Y(_08628_));
 sky130_fd_sc_hd__xnor2_1 _15534_ (.A(_08603_),
    .B(_08612_),
    .Y(_08629_));
 sky130_fd_sc_hd__and3_1 _15535_ (.A(_08599_),
    .B(_08592_),
    .C(_08598_),
    .X(_08630_));
 sky130_fd_sc_hd__a21oi_1 _15536_ (.A1(_08599_),
    .A2(_08592_),
    .B1(_08598_),
    .Y(_08631_));
 sky130_fd_sc_hd__or2_1 _15537_ (.A(_08630_),
    .B(_08631_),
    .X(_08632_));
 sky130_fd_sc_hd__and2b_1 _15538_ (.A_N(_08590_),
    .B(_08584_),
    .X(_08633_));
 sky130_fd_sc_hd__xnor2_1 _15539_ (.A(_08633_),
    .B(_08589_),
    .Y(_08634_));
 sky130_fd_sc_hd__xnor2_2 _15540_ (.A(_08578_),
    .B(_08579_),
    .Y(_08635_));
 sky130_fd_sc_hd__or4_1 _15541_ (.A(_08404_),
    .B(_08381_),
    .C(_08460_),
    .D(_08456_),
    .X(_08636_));
 sky130_fd_sc_hd__inv_2 _15542_ (.A(_08581_),
    .Y(_08637_));
 sky130_fd_sc_hd__a2bb2o_1 _15543_ (.A1_N(_08404_),
    .A2_N(_08472_),
    .B1(_08637_),
    .B2(_08380_),
    .X(_08638_));
 sky130_fd_sc_hd__or4bb_1 _15544_ (.A(_08178_),
    .B(_08439_),
    .C_N(_08636_),
    .D_N(_08638_),
    .X(_08639_));
 sky130_fd_sc_hd__and2_1 _15545_ (.A(_08636_),
    .B(_08639_),
    .X(_08640_));
 sky130_fd_sc_hd__xor2_1 _15546_ (.A(_08635_),
    .B(_08640_),
    .X(_08641_));
 sky130_fd_sc_hd__nand2_1 _15547_ (.A(_08237_),
    .B(_08214_),
    .Y(_08642_));
 sky130_fd_sc_hd__xnor2_1 _15548_ (.A(_08642_),
    .B(_08236_),
    .Y(_08643_));
 sky130_fd_sc_hd__nor2_1 _15549_ (.A(_08635_),
    .B(_08640_),
    .Y(_08644_));
 sky130_fd_sc_hd__a21oi_1 _15550_ (.A1(_08641_),
    .A2(_08643_),
    .B1(_08644_),
    .Y(_08645_));
 sky130_fd_sc_hd__xor2_1 _15551_ (.A(_08634_),
    .B(_08645_),
    .X(_08646_));
 sky130_fd_sc_hd__xnor2_1 _15552_ (.A(_08301_),
    .B(_08290_),
    .Y(_08647_));
 sky130_fd_sc_hd__nor2_1 _15553_ (.A(_08634_),
    .B(_08645_),
    .Y(_08648_));
 sky130_fd_sc_hd__a21oi_1 _15554_ (.A1(_08646_),
    .A2(_08647_),
    .B1(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__xor2_1 _15555_ (.A(_08632_),
    .B(_08649_),
    .X(_08650_));
 sky130_fd_sc_hd__xnor2_1 _15556_ (.A(_08364_),
    .B(_08354_),
    .Y(_08651_));
 sky130_fd_sc_hd__nand2_1 _15557_ (.A(_08650_),
    .B(_08651_),
    .Y(_08652_));
 sky130_fd_sc_hd__o21a_1 _15558_ (.A1(_08632_),
    .A2(_08649_),
    .B1(_08652_),
    .X(_08653_));
 sky130_fd_sc_hd__xor2_1 _15559_ (.A(_08629_),
    .B(_08653_),
    .X(_08654_));
 sky130_fd_sc_hd__nand2_1 _15560_ (.A(_08172_),
    .B(_08366_),
    .Y(_08655_));
 sky130_fd_sc_hd__and2_1 _15561_ (.A(_08367_),
    .B(_08655_),
    .X(_08656_));
 sky130_fd_sc_hd__o2bb2a_1 _15562_ (.A1_N(_08654_),
    .A2_N(_08656_),
    .B1(_08629_),
    .B2(_08653_),
    .X(_08657_));
 sky130_fd_sc_hd__xor2_1 _15563_ (.A(_08628_),
    .B(_08657_),
    .X(_08658_));
 sky130_fd_sc_hd__xnor2_2 _15564_ (.A(_08367_),
    .B(_08658_),
    .Y(_08659_));
 sky130_fd_sc_hd__or2_1 _15565_ (.A(_08650_),
    .B(_08651_),
    .X(_08660_));
 sky130_fd_sc_hd__nand2_1 _15566_ (.A(_08652_),
    .B(_08660_),
    .Y(_08661_));
 sky130_fd_sc_hd__xnor2_1 _15567_ (.A(_08646_),
    .B(_08647_),
    .Y(_08662_));
 sky130_fd_sc_hd__xnor2_1 _15568_ (.A(_08641_),
    .B(_08643_),
    .Y(_08663_));
 sky130_fd_sc_hd__a2bb2o_1 _15569_ (.A1_N(_08178_),
    .A2_N(_08440_),
    .B1(_08636_),
    .B2(_08638_),
    .X(_08664_));
 sky130_fd_sc_hd__or4_1 _15570_ (.A(_08177_),
    .B(_08382_),
    .C(_08461_),
    .D(_08457_),
    .X(_08665_));
 sky130_fd_sc_hd__clkbuf_4 _15571_ (.A(_08177_),
    .X(_08666_));
 sky130_fd_sc_hd__o22ai_1 _15572_ (.A1(_08382_),
    .A2(_08461_),
    .B1(_08457_),
    .B2(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__or4bb_1 _15573_ (.A(_08201_),
    .B(_08439_),
    .C_N(_08665_),
    .D_N(_08667_),
    .X(_08668_));
 sky130_fd_sc_hd__nand2_1 _15574_ (.A(_08665_),
    .B(_08668_),
    .Y(_08669_));
 sky130_fd_sc_hd__nand3_1 _15575_ (.A(_08639_),
    .B(_08664_),
    .C(_08669_),
    .Y(_08670_));
 sky130_fd_sc_hd__or2_1 _15576_ (.A(_08227_),
    .B(_08252_),
    .X(_08671_));
 sky130_fd_sc_hd__or3_1 _15577_ (.A(_08194_),
    .B(_08229_),
    .C(_08233_),
    .X(_08672_));
 sky130_fd_sc_hd__or3_1 _15578_ (.A(_08212_),
    .B(_08201_),
    .C(_08672_),
    .X(_08673_));
 sky130_fd_sc_hd__o22ai_1 _15579_ (.A1(_08195_),
    .A2(_08201_),
    .B1(_08234_),
    .B2(_08213_),
    .Y(_08674_));
 sky130_fd_sc_hd__and2_1 _15580_ (.A(_08673_),
    .B(_08674_),
    .X(_08675_));
 sky130_fd_sc_hd__xnor2_1 _15581_ (.A(_08671_),
    .B(_08675_),
    .Y(_08676_));
 sky130_fd_sc_hd__a21o_1 _15582_ (.A1(_08639_),
    .A2(_08664_),
    .B1(_08669_),
    .X(_08677_));
 sky130_fd_sc_hd__nand3_1 _15583_ (.A(_08670_),
    .B(_08676_),
    .C(_08677_),
    .Y(_08678_));
 sky130_fd_sc_hd__and2_1 _15584_ (.A(_08670_),
    .B(_08678_),
    .X(_08679_));
 sky130_fd_sc_hd__xor2_1 _15585_ (.A(_08663_),
    .B(_08679_),
    .X(_08680_));
 sky130_fd_sc_hd__nor2_1 _15586_ (.A(_08245_),
    .B(_08275_),
    .Y(_08681_));
 sky130_fd_sc_hd__nor2_1 _15587_ (.A(_08265_),
    .B(_08298_),
    .Y(_08682_));
 sky130_fd_sc_hd__nor2_1 _15588_ (.A(_08287_),
    .B(_08336_),
    .Y(_08683_));
 sky130_fd_sc_hd__xor2_1 _15589_ (.A(_08681_),
    .B(_08682_),
    .X(_08684_));
 sky130_fd_sc_hd__a22o_1 _15590_ (.A1(_08681_),
    .A2(_08682_),
    .B1(_08683_),
    .B2(_08684_),
    .X(_08685_));
 sky130_fd_sc_hd__or2b_1 _15591_ (.A(_08671_),
    .B_N(_08675_),
    .X(_08686_));
 sky130_fd_sc_hd__nand2_1 _15592_ (.A(_08300_),
    .B(_08291_),
    .Y(_08687_));
 sky130_fd_sc_hd__xor2_1 _15593_ (.A(_08687_),
    .B(_08299_),
    .X(_08688_));
 sky130_fd_sc_hd__a21o_1 _15594_ (.A1(_08673_),
    .A2(_08686_),
    .B1(_08688_),
    .X(_08689_));
 sky130_fd_sc_hd__nand3_1 _15595_ (.A(_08673_),
    .B(_08686_),
    .C(_08688_),
    .Y(_08690_));
 sky130_fd_sc_hd__nand2_1 _15596_ (.A(_08689_),
    .B(_08690_),
    .Y(_08691_));
 sky130_fd_sc_hd__xnor2_1 _15597_ (.A(_08685_),
    .B(_08691_),
    .Y(_08692_));
 sky130_fd_sc_hd__nor2_1 _15598_ (.A(_08663_),
    .B(_08679_),
    .Y(_08693_));
 sky130_fd_sc_hd__a21oi_1 _15599_ (.A1(_08680_),
    .A2(_08692_),
    .B1(_08693_),
    .Y(_08694_));
 sky130_fd_sc_hd__xor2_1 _15600_ (.A(_08662_),
    .B(_08694_),
    .X(_08695_));
 sky130_fd_sc_hd__buf_2 _15601_ (.A(_08358_),
    .X(_08696_));
 sky130_fd_sc_hd__nor2_1 _15602_ (.A(_08327_),
    .B(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__a21oi_1 _15603_ (.A1(_08346_),
    .A2(_08356_),
    .B1(_08360_),
    .Y(_08698_));
 sky130_fd_sc_hd__xnor2_1 _15604_ (.A(_08359_),
    .B(_08698_),
    .Y(_08699_));
 sky130_fd_sc_hd__and3_1 _15605_ (.A(_08356_),
    .B(_08697_),
    .C(_08699_),
    .X(_08700_));
 sky130_fd_sc_hd__a21bo_1 _15606_ (.A1(_08685_),
    .A2(_08690_),
    .B1_N(_08689_),
    .X(_08701_));
 sky130_fd_sc_hd__o21ai_2 _15607_ (.A1(_08152_),
    .A2(_08616_),
    .B1(_08362_),
    .Y(_08702_));
 sky130_fd_sc_hd__nand2_1 _15608_ (.A(_08363_),
    .B(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__xnor2_2 _15609_ (.A(_08701_),
    .B(_08703_),
    .Y(_08704_));
 sky130_fd_sc_hd__xor2_1 _15610_ (.A(_08700_),
    .B(_08704_),
    .X(_08705_));
 sky130_fd_sc_hd__nor2_1 _15611_ (.A(_08662_),
    .B(_08694_),
    .Y(_08706_));
 sky130_fd_sc_hd__a21oi_1 _15612_ (.A1(_08695_),
    .A2(_08705_),
    .B1(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__xnor2_2 _15613_ (.A(_08661_),
    .B(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__a32oi_4 _15614_ (.A1(_08363_),
    .A2(_08701_),
    .A3(_08702_),
    .B1(_08704_),
    .B2(_08700_),
    .Y(_08709_));
 sky130_fd_sc_hd__xnor2_2 _15615_ (.A(_08708_),
    .B(_08709_),
    .Y(_08710_));
 sky130_fd_sc_hd__xnor2_1 _15616_ (.A(_08683_),
    .B(_08684_),
    .Y(_08711_));
 sky130_fd_sc_hd__or3b_1 _15617_ (.A(_08213_),
    .B(_08250_),
    .C_N(_08251_),
    .X(_08712_));
 sky130_fd_sc_hd__xor2_1 _15618_ (.A(_08672_),
    .B(_08712_),
    .X(_08713_));
 sky130_fd_sc_hd__nor2_1 _15619_ (.A(_08227_),
    .B(_08276_),
    .Y(_08714_));
 sky130_fd_sc_hd__a2bb2o_1 _15620_ (.A1_N(_08672_),
    .A2_N(_08712_),
    .B1(_08713_),
    .B2(_08714_),
    .X(_08715_));
 sky130_fd_sc_hd__or2b_1 _15621_ (.A(_08711_),
    .B_N(_08715_),
    .X(_08716_));
 sky130_fd_sc_hd__xor2_1 _15622_ (.A(_08715_),
    .B(_08711_),
    .X(_08717_));
 sky130_fd_sc_hd__a211o_1 _15623_ (.A1(_08292_),
    .A2(_08357_),
    .B1(_08245_),
    .C1(_08296_),
    .X(_08718_));
 sky130_fd_sc_hd__or3_2 _15624_ (.A(_08265_),
    .B(_08332_),
    .C(_08335_),
    .X(_08719_));
 sky130_fd_sc_hd__nor2_1 _15625_ (.A(_08287_),
    .B(_08343_),
    .Y(_08720_));
 sky130_fd_sc_hd__xor2_1 _15626_ (.A(_08718_),
    .B(_08719_),
    .X(_08721_));
 sky130_fd_sc_hd__a2bb2o_1 _15627_ (.A1_N(_08718_),
    .A2_N(_08719_),
    .B1(_08720_),
    .B2(_08721_),
    .X(_08722_));
 sky130_fd_sc_hd__or2b_1 _15628_ (.A(_08717_),
    .B_N(_08722_),
    .X(_08723_));
 sky130_fd_sc_hd__a21oi_1 _15629_ (.A1(_08356_),
    .A2(_08697_),
    .B1(_08699_),
    .Y(_08724_));
 sky130_fd_sc_hd__or2_1 _15630_ (.A(_08700_),
    .B(_08724_),
    .X(_08725_));
 sky130_fd_sc_hd__a21oi_2 _15631_ (.A1(_08716_),
    .A2(_08723_),
    .B1(_08725_),
    .Y(_08726_));
 sky130_fd_sc_hd__xnor2_1 _15632_ (.A(_08695_),
    .B(_08705_),
    .Y(_08727_));
 sky130_fd_sc_hd__xnor2_1 _15633_ (.A(_08680_),
    .B(_08692_),
    .Y(_08728_));
 sky130_fd_sc_hd__a21o_1 _15634_ (.A1(_08670_),
    .A2(_08677_),
    .B1(_08676_),
    .X(_08729_));
 sky130_fd_sc_hd__a2bb2o_1 _15635_ (.A1_N(_08201_),
    .A2_N(_08440_),
    .B1(_08665_),
    .B2(_08667_),
    .X(_08730_));
 sky130_fd_sc_hd__clkbuf_4 _15636_ (.A(_08233_),
    .X(_08731_));
 sky130_fd_sc_hd__nor2_1 _15637_ (.A(_08229_),
    .B(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__a221o_4 _15638_ (.A1(\rbzero.wall_tracer.visualWallDist[-9] ),
    .A2(_08149_),
    .B1(_08357_),
    .B2(\rbzero.debug_overlay.playerX[-9] ),
    .C1(_08438_),
    .X(_08733_));
 sky130_fd_sc_hd__clkbuf_4 _15639_ (.A(_08200_),
    .X(_08734_));
 sky130_fd_sc_hd__o22ai_2 _15640_ (.A1(_08666_),
    .A2(_08472_),
    .B1(_08457_),
    .B2(_08734_),
    .Y(_08735_));
 sky130_fd_sc_hd__and4bb_1 _15641_ (.A_N(_08666_),
    .B_N(_08734_),
    .C(_08484_),
    .D(_08471_),
    .X(_08736_));
 sky130_fd_sc_hd__a31o_1 _15642_ (.A1(_08732_),
    .A2(_08733_),
    .A3(_08735_),
    .B1(_08736_),
    .X(_08737_));
 sky130_fd_sc_hd__nand3_1 _15643_ (.A(_08668_),
    .B(_08730_),
    .C(_08737_),
    .Y(_08738_));
 sky130_fd_sc_hd__xor2_1 _15644_ (.A(_08714_),
    .B(_08713_),
    .X(_08739_));
 sky130_fd_sc_hd__a21o_1 _15645_ (.A1(_08668_),
    .A2(_08730_),
    .B1(_08737_),
    .X(_08740_));
 sky130_fd_sc_hd__nand3_1 _15646_ (.A(_08738_),
    .B(_08739_),
    .C(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__nand2_1 _15647_ (.A(_08738_),
    .B(_08741_),
    .Y(_08742_));
 sky130_fd_sc_hd__nand3_1 _15648_ (.A(_08678_),
    .B(_08729_),
    .C(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__xnor2_1 _15649_ (.A(_08722_),
    .B(_08717_),
    .Y(_08744_));
 sky130_fd_sc_hd__a21o_1 _15650_ (.A1(_08678_),
    .A2(_08729_),
    .B1(_08742_),
    .X(_08745_));
 sky130_fd_sc_hd__nand3_1 _15651_ (.A(_08743_),
    .B(_08744_),
    .C(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__and2_1 _15652_ (.A(_08743_),
    .B(_08746_),
    .X(_08747_));
 sky130_fd_sc_hd__xor2_1 _15653_ (.A(_08728_),
    .B(_08747_),
    .X(_08748_));
 sky130_fd_sc_hd__and3_1 _15654_ (.A(_08716_),
    .B(_08723_),
    .C(_08725_),
    .X(_08749_));
 sky130_fd_sc_hd__nor2_1 _15655_ (.A(_08726_),
    .B(_08749_),
    .Y(_08750_));
 sky130_fd_sc_hd__nor2_1 _15656_ (.A(_08728_),
    .B(_08747_),
    .Y(_08751_));
 sky130_fd_sc_hd__a21o_1 _15657_ (.A1(_08748_),
    .A2(_08750_),
    .B1(_08751_),
    .X(_08752_));
 sky130_fd_sc_hd__xnor2_1 _15658_ (.A(_08727_),
    .B(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__or2b_1 _15659_ (.A(_08727_),
    .B_N(_08752_),
    .X(_08754_));
 sky130_fd_sc_hd__a21boi_2 _15660_ (.A1(_08726_),
    .A2(_08753_),
    .B1_N(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__nor2_1 _15661_ (.A(_08710_),
    .B(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__inv_2 _15662_ (.A(_08756_),
    .Y(_08757_));
 sky130_fd_sc_hd__xnor2_1 _15663_ (.A(_08654_),
    .B(_08656_),
    .Y(_08758_));
 sky130_fd_sc_hd__or2_1 _15664_ (.A(_08661_),
    .B(_08707_),
    .X(_08759_));
 sky130_fd_sc_hd__o21a_1 _15665_ (.A1(_08708_),
    .A2(_08709_),
    .B1(_08759_),
    .X(_08760_));
 sky130_fd_sc_hd__nor2_1 _15666_ (.A(_08758_),
    .B(_08760_),
    .Y(_08761_));
 sky130_fd_sc_hd__and2_1 _15667_ (.A(_08758_),
    .B(_08760_),
    .X(_08762_));
 sky130_fd_sc_hd__or2_1 _15668_ (.A(_08761_),
    .B(_08762_),
    .X(_08763_));
 sky130_fd_sc_hd__nor2_1 _15669_ (.A(_08757_),
    .B(_08763_),
    .Y(_08764_));
 sky130_fd_sc_hd__xnor2_1 _15670_ (.A(_08726_),
    .B(_08753_),
    .Y(_08765_));
 sky130_fd_sc_hd__or2_1 _15671_ (.A(_08195_),
    .B(_08275_),
    .X(_08766_));
 sky130_fd_sc_hd__or3b_1 _15672_ (.A(_08195_),
    .B(_08250_),
    .C_N(_08251_),
    .X(_08767_));
 sky130_fd_sc_hd__or3_1 _15673_ (.A(_08213_),
    .B(_08269_),
    .C(_08274_),
    .X(_08768_));
 sky130_fd_sc_hd__xor2_1 _15674_ (.A(_08767_),
    .B(_08768_),
    .X(_08769_));
 sky130_fd_sc_hd__nor2_1 _15675_ (.A(_08228_),
    .B(_08298_),
    .Y(_08770_));
 sky130_fd_sc_hd__a2bb2oi_1 _15676_ (.A1_N(_08712_),
    .A2_N(_08766_),
    .B1(_08769_),
    .B2(_08770_),
    .Y(_08771_));
 sky130_fd_sc_hd__xnor2_1 _15677_ (.A(_08720_),
    .B(_08721_),
    .Y(_08772_));
 sky130_fd_sc_hd__or2_1 _15678_ (.A(_08771_),
    .B(_08772_),
    .X(_08773_));
 sky130_fd_sc_hd__o22a_1 _15679_ (.A1(_08246_),
    .A2(_08337_),
    .B1(_08343_),
    .B2(_08265_),
    .X(_08774_));
 sky130_fd_sc_hd__or3_1 _15680_ (.A(_08246_),
    .B(_08343_),
    .C(_08719_),
    .X(_08775_));
 sky130_fd_sc_hd__o31a_1 _15681_ (.A1(_08287_),
    .A2(_08358_),
    .A3(_08774_),
    .B1(_08775_),
    .X(_08776_));
 sky130_fd_sc_hd__xnor2_1 _15682_ (.A(_08771_),
    .B(_08772_),
    .Y(_08777_));
 sky130_fd_sc_hd__or2_1 _15683_ (.A(_08776_),
    .B(_08777_),
    .X(_08778_));
 sky130_fd_sc_hd__nand2_1 _15684_ (.A(_08356_),
    .B(_08697_),
    .Y(_08779_));
 sky130_fd_sc_hd__or2_1 _15685_ (.A(_08356_),
    .B(_08697_),
    .X(_08780_));
 sky130_fd_sc_hd__nand2_1 _15686_ (.A(_08779_),
    .B(_08780_),
    .Y(_08781_));
 sky130_fd_sc_hd__a21oi_2 _15687_ (.A1(_08773_),
    .A2(_08778_),
    .B1(_08781_),
    .Y(_08782_));
 sky130_fd_sc_hd__xnor2_1 _15688_ (.A(_08748_),
    .B(_08750_),
    .Y(_08783_));
 sky130_fd_sc_hd__a21o_1 _15689_ (.A1(_08743_),
    .A2(_08745_),
    .B1(_08744_),
    .X(_08784_));
 sky130_fd_sc_hd__a21o_1 _15690_ (.A1(_08738_),
    .A2(_08740_),
    .B1(_08739_),
    .X(_08785_));
 sky130_fd_sc_hd__xor2_1 _15691_ (.A(_08770_),
    .B(_08769_),
    .X(_08786_));
 sky130_fd_sc_hd__or4b_1 _15692_ (.A(_08235_),
    .B(_08440_),
    .C(_08736_),
    .D_N(_08735_),
    .X(_08787_));
 sky130_fd_sc_hd__or4_1 _15693_ (.A(_08666_),
    .B(_08734_),
    .C(_08472_),
    .D(_08457_),
    .X(_08788_));
 sky130_fd_sc_hd__a22o_1 _15694_ (.A1(_08732_),
    .A2(_08733_),
    .B1(_08788_),
    .B2(_08735_),
    .X(_08789_));
 sky130_fd_sc_hd__o22ai_2 _15695_ (.A1(_08734_),
    .A2(_08473_),
    .B1(_08457_),
    .B2(_08233_),
    .Y(_08790_));
 sky130_fd_sc_hd__and4bb_1 _15696_ (.A_N(_08734_),
    .B_N(_08233_),
    .C(_08484_),
    .D(_08471_),
    .X(_08791_));
 sky130_fd_sc_hd__a31o_1 _15697_ (.A1(_08529_),
    .A2(_08733_),
    .A3(_08790_),
    .B1(_08791_),
    .X(_08792_));
 sky130_fd_sc_hd__a21o_1 _15698_ (.A1(_08787_),
    .A2(_08789_),
    .B1(_08792_),
    .X(_08793_));
 sky130_fd_sc_hd__and3_1 _15699_ (.A(_08787_),
    .B(_08789_),
    .C(_08792_),
    .X(_08794_));
 sky130_fd_sc_hd__a21o_1 _15700_ (.A1(_08786_),
    .A2(_08793_),
    .B1(_08794_),
    .X(_08795_));
 sky130_fd_sc_hd__nand3_1 _15701_ (.A(_08741_),
    .B(_08785_),
    .C(_08795_),
    .Y(_08796_));
 sky130_fd_sc_hd__xor2_1 _15702_ (.A(_08776_),
    .B(_08777_),
    .X(_08797_));
 sky130_fd_sc_hd__a21o_1 _15703_ (.A1(_08741_),
    .A2(_08785_),
    .B1(_08795_),
    .X(_08798_));
 sky130_fd_sc_hd__nand3_1 _15704_ (.A(_08796_),
    .B(_08797_),
    .C(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__nand2_1 _15705_ (.A(_08796_),
    .B(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__a21o_1 _15706_ (.A1(_08746_),
    .A2(_08784_),
    .B1(_08800_),
    .X(_08801_));
 sky130_fd_sc_hd__and3_1 _15707_ (.A(_08773_),
    .B(_08778_),
    .C(_08781_),
    .X(_08802_));
 sky130_fd_sc_hd__nor2_1 _15708_ (.A(_08782_),
    .B(_08802_),
    .Y(_08803_));
 sky130_fd_sc_hd__nand3_1 _15709_ (.A(_08746_),
    .B(_08784_),
    .C(_08800_),
    .Y(_08804_));
 sky130_fd_sc_hd__a21boi_1 _15710_ (.A1(_08801_),
    .A2(_08803_),
    .B1_N(_08804_),
    .Y(_08805_));
 sky130_fd_sc_hd__xor2_1 _15711_ (.A(_08783_),
    .B(_08805_),
    .X(_08806_));
 sky130_fd_sc_hd__nor2_1 _15712_ (.A(_08783_),
    .B(_08805_),
    .Y(_08807_));
 sky130_fd_sc_hd__a21oi_1 _15713_ (.A1(_08782_),
    .A2(_08806_),
    .B1(_08807_),
    .Y(_08808_));
 sky130_fd_sc_hd__nor2_1 _15714_ (.A(_08765_),
    .B(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__xor2_2 _15715_ (.A(_08710_),
    .B(_08755_),
    .X(_08810_));
 sky130_fd_sc_hd__nand2_1 _15716_ (.A(_08809_),
    .B(_08810_),
    .Y(_08811_));
 sky130_fd_sc_hd__xnor2_1 _15717_ (.A(_08782_),
    .B(_08806_),
    .Y(_08812_));
 sky130_fd_sc_hd__clkbuf_4 _15718_ (.A(_08328_),
    .X(_08813_));
 sky130_fd_sc_hd__buf_4 _15719_ (.A(_08813_),
    .X(_08814_));
 sky130_fd_sc_hd__or2_1 _15720_ (.A(_08814_),
    .B(_08696_),
    .X(_08815_));
 sky130_fd_sc_hd__clkbuf_4 _15721_ (.A(_08516_),
    .X(_08816_));
 sky130_fd_sc_hd__or2_1 _15722_ (.A(_08213_),
    .B(_08297_),
    .X(_08817_));
 sky130_fd_sc_hd__or2_1 _15723_ (.A(_08228_),
    .B(_08336_),
    .X(_08818_));
 sky130_fd_sc_hd__xor2_1 _15724_ (.A(_08766_),
    .B(_08817_),
    .X(_08819_));
 sky130_fd_sc_hd__or2b_1 _15725_ (.A(_08818_),
    .B_N(_08819_),
    .X(_08820_));
 sky130_fd_sc_hd__o21a_1 _15726_ (.A1(_08766_),
    .A2(_08817_),
    .B1(_08820_),
    .X(_08821_));
 sky130_fd_sc_hd__or2_1 _15727_ (.A(_08287_),
    .B(_08358_),
    .X(_08822_));
 sky130_fd_sc_hd__nor3_1 _15728_ (.A(_08246_),
    .B(_08344_),
    .C(_08719_),
    .Y(_08823_));
 sky130_fd_sc_hd__nor2_1 _15729_ (.A(_08823_),
    .B(_08774_),
    .Y(_08824_));
 sky130_fd_sc_hd__xnor2_1 _15730_ (.A(_08822_),
    .B(_08824_),
    .Y(_08825_));
 sky130_fd_sc_hd__xor2_1 _15731_ (.A(_08821_),
    .B(_08825_),
    .X(_08826_));
 sky130_fd_sc_hd__or2_1 _15732_ (.A(_08369_),
    .B(_08696_),
    .X(_08827_));
 sky130_fd_sc_hd__or2b_1 _15733_ (.A(_08821_),
    .B_N(_08825_),
    .X(_08828_));
 sky130_fd_sc_hd__o41a_1 _15734_ (.A1(_08816_),
    .A2(_08344_),
    .A3(_08826_),
    .A4(_08827_),
    .B1(_08828_),
    .X(_08829_));
 sky130_fd_sc_hd__nor2_1 _15735_ (.A(_08815_),
    .B(_08829_),
    .Y(_08830_));
 sky130_fd_sc_hd__and3_1 _15736_ (.A(_08804_),
    .B(_08801_),
    .C(_08803_),
    .X(_08831_));
 sky130_fd_sc_hd__a21oi_1 _15737_ (.A1(_08804_),
    .A2(_08801_),
    .B1(_08803_),
    .Y(_08832_));
 sky130_fd_sc_hd__or2_1 _15738_ (.A(_08831_),
    .B(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__and2_1 _15739_ (.A(_08815_),
    .B(_08829_),
    .X(_08834_));
 sky130_fd_sc_hd__nor2_1 _15740_ (.A(_08830_),
    .B(_08834_),
    .Y(_08835_));
 sky130_fd_sc_hd__a21o_1 _15741_ (.A1(_08796_),
    .A2(_08798_),
    .B1(_08797_),
    .X(_08836_));
 sky130_fd_sc_hd__nand2_1 _15742_ (.A(_08799_),
    .B(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__nor3_1 _15743_ (.A(_08516_),
    .B(_08344_),
    .C(_08827_),
    .Y(_08838_));
 sky130_fd_sc_hd__xnor2_1 _15744_ (.A(_08826_),
    .B(_08838_),
    .Y(_08839_));
 sky130_fd_sc_hd__inv_2 _15745_ (.A(_08794_),
    .Y(_08840_));
 sky130_fd_sc_hd__nand3_1 _15746_ (.A(_08840_),
    .B(_08786_),
    .C(_08793_),
    .Y(_08841_));
 sky130_fd_sc_hd__a21o_1 _15747_ (.A1(_08840_),
    .A2(_08793_),
    .B1(_08786_),
    .X(_08842_));
 sky130_fd_sc_hd__or4b_1 _15748_ (.A(_08252_),
    .B(_08440_),
    .C(_08791_),
    .D_N(_08790_),
    .X(_08843_));
 sky130_fd_sc_hd__or4_1 _15749_ (.A(_08734_),
    .B(_08233_),
    .C(_08472_),
    .D(_08457_),
    .X(_08844_));
 sky130_fd_sc_hd__a22o_1 _15750_ (.A1(_08529_),
    .A2(_08733_),
    .B1(_08844_),
    .B2(_08790_),
    .X(_08845_));
 sky130_fd_sc_hd__nor2_1 _15751_ (.A(_08276_),
    .B(_08440_),
    .Y(_08846_));
 sky130_fd_sc_hd__clkbuf_4 _15752_ (.A(_08250_),
    .X(_08847_));
 sky130_fd_sc_hd__o22ai_1 _15753_ (.A1(_08731_),
    .A2(_08473_),
    .B1(_08457_),
    .B2(_08847_),
    .Y(_08848_));
 sky130_fd_sc_hd__or4_1 _15754_ (.A(_08731_),
    .B(_08847_),
    .C(_08473_),
    .D(_08457_),
    .X(_08849_));
 sky130_fd_sc_hd__a21bo_1 _15755_ (.A1(_08846_),
    .A2(_08848_),
    .B1_N(_08849_),
    .X(_08850_));
 sky130_fd_sc_hd__xnor2_1 _15756_ (.A(_08818_),
    .B(_08819_),
    .Y(_08851_));
 sky130_fd_sc_hd__nand2_1 _15757_ (.A(_08843_),
    .B(_08845_),
    .Y(_08852_));
 sky130_fd_sc_hd__xnor2_1 _15758_ (.A(_08852_),
    .B(_08850_),
    .Y(_08853_));
 sky130_fd_sc_hd__a32o_1 _15759_ (.A1(_08843_),
    .A2(_08845_),
    .A3(_08850_),
    .B1(_08851_),
    .B2(_08853_),
    .X(_08854_));
 sky130_fd_sc_hd__a21o_1 _15760_ (.A1(_08841_),
    .A2(_08842_),
    .B1(_08854_),
    .X(_08855_));
 sky130_fd_sc_hd__and3_1 _15761_ (.A(_08841_),
    .B(_08842_),
    .C(_08854_),
    .X(_08856_));
 sky130_fd_sc_hd__a21o_1 _15762_ (.A1(_08839_),
    .A2(_08855_),
    .B1(_08856_),
    .X(_08857_));
 sky130_fd_sc_hd__xnor2_1 _15763_ (.A(_08837_),
    .B(_08857_),
    .Y(_08858_));
 sky130_fd_sc_hd__and3_1 _15764_ (.A(_08799_),
    .B(_08836_),
    .C(_08857_),
    .X(_08859_));
 sky130_fd_sc_hd__a21oi_1 _15765_ (.A1(_08835_),
    .A2(_08858_),
    .B1(_08859_),
    .Y(_08860_));
 sky130_fd_sc_hd__xor2_1 _15766_ (.A(_08833_),
    .B(_08860_),
    .X(_08861_));
 sky130_fd_sc_hd__nor2_1 _15767_ (.A(_08833_),
    .B(_08860_),
    .Y(_08862_));
 sky130_fd_sc_hd__a21oi_1 _15768_ (.A1(_08830_),
    .A2(_08861_),
    .B1(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__nor2_1 _15769_ (.A(_08812_),
    .B(_08863_),
    .Y(_08864_));
 sky130_fd_sc_hd__xor2_1 _15770_ (.A(_08765_),
    .B(_08808_),
    .X(_08865_));
 sky130_fd_sc_hd__and2_1 _15771_ (.A(_08864_),
    .B(_08865_),
    .X(_08866_));
 sky130_fd_sc_hd__xor2_1 _15772_ (.A(_08812_),
    .B(_08863_),
    .X(_08867_));
 sky130_fd_sc_hd__xor2_1 _15773_ (.A(_08830_),
    .B(_08861_),
    .X(_08868_));
 sky130_fd_sc_hd__or2b_1 _15774_ (.A(_08856_),
    .B_N(_08855_),
    .X(_08869_));
 sky130_fd_sc_hd__xor2_1 _15775_ (.A(_08839_),
    .B(_08869_),
    .X(_08870_));
 sky130_fd_sc_hd__xnor2_1 _15776_ (.A(_08851_),
    .B(_08853_),
    .Y(_08871_));
 sky130_fd_sc_hd__nand2_1 _15777_ (.A(_08849_),
    .B(_08848_),
    .Y(_08872_));
 sky130_fd_sc_hd__xor2_1 _15778_ (.A(_08846_),
    .B(_08872_),
    .X(_08873_));
 sky130_fd_sc_hd__nor2_1 _15779_ (.A(_08298_),
    .B(_08441_),
    .Y(_08874_));
 sky130_fd_sc_hd__nor4_1 _15780_ (.A(_08039_),
    .B(_08847_),
    .C(_08274_),
    .D(_08458_),
    .Y(_08875_));
 sky130_fd_sc_hd__o22a_1 _15781_ (.A1(_08847_),
    .A2(_08473_),
    .B1(_08458_),
    .B2(_08274_),
    .X(_08876_));
 sky130_fd_sc_hd__nor2_1 _15782_ (.A(_08875_),
    .B(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__a21oi_1 _15783_ (.A1(_08874_),
    .A2(_08877_),
    .B1(_08875_),
    .Y(_08878_));
 sky130_fd_sc_hd__xor2_1 _15784_ (.A(_08873_),
    .B(_08878_),
    .X(_08879_));
 sky130_fd_sc_hd__or2_1 _15785_ (.A(_08228_),
    .B(_08344_),
    .X(_08880_));
 sky130_fd_sc_hd__o22a_1 _15786_ (.A1(_08195_),
    .A2(_08298_),
    .B1(_08337_),
    .B2(_08410_),
    .X(_08881_));
 sky130_fd_sc_hd__or4_1 _15787_ (.A(_08213_),
    .B(_08195_),
    .C(_08298_),
    .D(_08337_),
    .X(_08882_));
 sky130_fd_sc_hd__and2b_1 _15788_ (.A_N(_08881_),
    .B(_08882_),
    .X(_08883_));
 sky130_fd_sc_hd__xnor2_1 _15789_ (.A(_08880_),
    .B(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__nand2_1 _15790_ (.A(_08879_),
    .B(_08884_),
    .Y(_08885_));
 sky130_fd_sc_hd__o21ai_1 _15791_ (.A1(_08873_),
    .A2(_08878_),
    .B1(_08885_),
    .Y(_08886_));
 sky130_fd_sc_hd__xnor2_1 _15792_ (.A(_08871_),
    .B(_08886_),
    .Y(_08887_));
 sky130_fd_sc_hd__o21ai_1 _15793_ (.A1(_08880_),
    .A2(_08881_),
    .B1(_08882_),
    .Y(_08888_));
 sky130_fd_sc_hd__buf_4 _15794_ (.A(_08369_),
    .X(_08889_));
 sky130_fd_sc_hd__o22a_1 _15795_ (.A1(_08889_),
    .A2(_08344_),
    .B1(_08696_),
    .B2(_08516_),
    .X(_08890_));
 sky130_fd_sc_hd__or2_1 _15796_ (.A(_08838_),
    .B(_08890_),
    .X(_08891_));
 sky130_fd_sc_hd__xnor2_1 _15797_ (.A(_08888_),
    .B(_08891_),
    .Y(_08892_));
 sky130_fd_sc_hd__and2b_1 _15798_ (.A_N(_08871_),
    .B(_08886_),
    .X(_08893_));
 sky130_fd_sc_hd__a21oi_1 _15799_ (.A1(_08887_),
    .A2(_08892_),
    .B1(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__or2_1 _15800_ (.A(_08870_),
    .B(_08894_),
    .X(_08895_));
 sky130_fd_sc_hd__and2b_1 _15801_ (.A_N(_08891_),
    .B(_08888_),
    .X(_08896_));
 sky130_fd_sc_hd__xor2_1 _15802_ (.A(_08870_),
    .B(_08894_),
    .X(_08897_));
 sky130_fd_sc_hd__nand2_1 _15803_ (.A(_08896_),
    .B(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__xnor2_1 _15804_ (.A(_08835_),
    .B(_08858_),
    .Y(_08899_));
 sky130_fd_sc_hd__a21o_1 _15805_ (.A1(_08895_),
    .A2(_08898_),
    .B1(_08899_),
    .X(_08900_));
 sky130_fd_sc_hd__inv_2 _15806_ (.A(_08900_),
    .Y(_08901_));
 sky130_fd_sc_hd__and2_1 _15807_ (.A(_08868_),
    .B(_08901_),
    .X(_08902_));
 sky130_fd_sc_hd__and2_1 _15808_ (.A(_08867_),
    .B(_08902_),
    .X(_08903_));
 sky130_fd_sc_hd__nor2_1 _15809_ (.A(_08864_),
    .B(_08903_),
    .Y(_08904_));
 sky130_fd_sc_hd__xnor2_1 _15810_ (.A(_08865_),
    .B(_08904_),
    .Y(_08905_));
 sky130_fd_sc_hd__xnor2_1 _15811_ (.A(_08867_),
    .B(_08902_),
    .Y(_08906_));
 sky130_fd_sc_hd__nand2_1 _15812_ (.A(_08899_),
    .B(_08895_),
    .Y(_08907_));
 sky130_fd_sc_hd__or2_1 _15813_ (.A(_08896_),
    .B(_08897_),
    .X(_08908_));
 sky130_fd_sc_hd__nand2_1 _15814_ (.A(_08898_),
    .B(_08908_),
    .Y(_08909_));
 sky130_fd_sc_hd__clkbuf_4 _15815_ (.A(_08410_),
    .X(_08910_));
 sky130_fd_sc_hd__or2_1 _15816_ (.A(_08195_),
    .B(_08337_),
    .X(_08911_));
 sky130_fd_sc_hd__nor2_1 _15817_ (.A(_08213_),
    .B(_08343_),
    .Y(_08912_));
 sky130_fd_sc_hd__xnor2_1 _15818_ (.A(_08911_),
    .B(_08912_),
    .Y(_08913_));
 sky130_fd_sc_hd__or3b_1 _15819_ (.A(_08228_),
    .B(_08696_),
    .C_N(_08913_),
    .X(_08914_));
 sky130_fd_sc_hd__o31a_1 _15820_ (.A1(_08910_),
    .A2(_08344_),
    .A3(_08911_),
    .B1(_08914_),
    .X(_08915_));
 sky130_fd_sc_hd__nor2_1 _15821_ (.A(_08827_),
    .B(_08915_),
    .Y(_08916_));
 sky130_fd_sc_hd__xnor2_1 _15822_ (.A(_08887_),
    .B(_08892_),
    .Y(_08917_));
 sky130_fd_sc_hd__or2_1 _15823_ (.A(_08879_),
    .B(_08884_),
    .X(_08918_));
 sky130_fd_sc_hd__nand2_1 _15824_ (.A(_08885_),
    .B(_08918_),
    .Y(_08919_));
 sky130_fd_sc_hd__xnor2_1 _15825_ (.A(_08874_),
    .B(_08877_),
    .Y(_08920_));
 sky130_fd_sc_hd__nor2_1 _15826_ (.A(_08337_),
    .B(_08441_),
    .Y(_08921_));
 sky130_fd_sc_hd__or4_1 _15827_ (.A(_08039_),
    .B(_08274_),
    .C(_08296_),
    .D(_08458_),
    .X(_08922_));
 sky130_fd_sc_hd__inv_2 _15828_ (.A(_08922_),
    .Y(_08923_));
 sky130_fd_sc_hd__o22a_1 _15829_ (.A1(_08274_),
    .A2(_08473_),
    .B1(_08458_),
    .B2(_08296_),
    .X(_08924_));
 sky130_fd_sc_hd__nor2_1 _15830_ (.A(_08923_),
    .B(_08924_),
    .Y(_08925_));
 sky130_fd_sc_hd__a21oi_1 _15831_ (.A1(_08921_),
    .A2(_08925_),
    .B1(_08923_),
    .Y(_08926_));
 sky130_fd_sc_hd__o21bai_1 _15832_ (.A1(_08434_),
    .A2(_08696_),
    .B1_N(_08913_),
    .Y(_08927_));
 sky130_fd_sc_hd__and2_1 _15833_ (.A(_08914_),
    .B(_08927_),
    .X(_08928_));
 sky130_fd_sc_hd__xor2_1 _15834_ (.A(_08920_),
    .B(_08926_),
    .X(_08929_));
 sky130_fd_sc_hd__nand2_1 _15835_ (.A(_08928_),
    .B(_08929_),
    .Y(_08930_));
 sky130_fd_sc_hd__o21a_1 _15836_ (.A1(_08920_),
    .A2(_08926_),
    .B1(_08930_),
    .X(_08931_));
 sky130_fd_sc_hd__xor2_1 _15837_ (.A(_08919_),
    .B(_08931_),
    .X(_08932_));
 sky130_fd_sc_hd__and2_1 _15838_ (.A(_08827_),
    .B(_08915_),
    .X(_08933_));
 sky130_fd_sc_hd__nor2_1 _15839_ (.A(_08916_),
    .B(_08933_),
    .Y(_08934_));
 sky130_fd_sc_hd__nand2_1 _15840_ (.A(_08932_),
    .B(_08934_),
    .Y(_08935_));
 sky130_fd_sc_hd__o21a_1 _15841_ (.A1(_08919_),
    .A2(_08931_),
    .B1(_08935_),
    .X(_08936_));
 sky130_fd_sc_hd__xor2_1 _15842_ (.A(_08917_),
    .B(_08936_),
    .X(_08937_));
 sky130_fd_sc_hd__or2_1 _15843_ (.A(_08917_),
    .B(_08936_),
    .X(_08938_));
 sky130_fd_sc_hd__a21boi_1 _15844_ (.A1(_08916_),
    .A2(_08937_),
    .B1_N(_08938_),
    .Y(_08939_));
 sky130_fd_sc_hd__nor2_1 _15845_ (.A(_08909_),
    .B(_08939_),
    .Y(_08940_));
 sky130_fd_sc_hd__and4_1 _15846_ (.A(_08868_),
    .B(_08900_),
    .C(_08907_),
    .D(_08940_),
    .X(_08941_));
 sky130_fd_sc_hd__xnor2_1 _15847_ (.A(_08906_),
    .B(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__nor2_1 _15848_ (.A(_08431_),
    .B(_08696_),
    .Y(_08943_));
 sky130_fd_sc_hd__nor2_1 _15849_ (.A(_08335_),
    .B(_08473_),
    .Y(_08944_));
 sky130_fd_sc_hd__nor2_1 _15850_ (.A(_08304_),
    .B(_08458_),
    .Y(_08945_));
 sky130_fd_sc_hd__xor2_1 _15851_ (.A(_08944_),
    .B(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__and3b_1 _15852_ (.A_N(_08696_),
    .B(_08733_),
    .C(_08946_),
    .X(_08947_));
 sky130_fd_sc_hd__a21o_1 _15853_ (.A1(_08944_),
    .A2(_08945_),
    .B1(_08947_),
    .X(_08948_));
 sky130_fd_sc_hd__nand2_1 _15854_ (.A(_08943_),
    .B(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__clkbuf_4 _15855_ (.A(_08441_),
    .X(_08950_));
 sky130_fd_sc_hd__nor2_1 _15856_ (.A(_08344_),
    .B(_08950_),
    .Y(_08951_));
 sky130_fd_sc_hd__buf_4 _15857_ (.A(_08296_),
    .X(_08952_));
 sky130_fd_sc_hd__nand2_1 _15858_ (.A(_08471_),
    .B(_08944_),
    .Y(_08953_));
 sky130_fd_sc_hd__o22a_1 _15859_ (.A1(_08296_),
    .A2(_08473_),
    .B1(_08458_),
    .B2(_08335_),
    .X(_08954_));
 sky130_fd_sc_hd__o21ba_1 _15860_ (.A1(_08952_),
    .A2(_08953_),
    .B1_N(_08954_),
    .X(_08955_));
 sky130_fd_sc_hd__xnor2_1 _15861_ (.A(_08951_),
    .B(_08955_),
    .Y(_08956_));
 sky130_fd_sc_hd__or3b_1 _15862_ (.A(_08616_),
    .B(_08461_),
    .C_N(_08945_),
    .X(_08957_));
 sky130_fd_sc_hd__o21ba_1 _15863_ (.A1(_08696_),
    .A2(_08950_),
    .B1_N(_08946_),
    .X(_08958_));
 sky130_fd_sc_hd__or3_1 _15864_ (.A(_08947_),
    .B(_08957_),
    .C(_08958_),
    .X(_08959_));
 sky130_fd_sc_hd__xnor2_1 _15865_ (.A(_08921_),
    .B(_08925_),
    .Y(_08960_));
 sky130_fd_sc_hd__or2_1 _15866_ (.A(_08296_),
    .B(_08953_),
    .X(_08961_));
 sky130_fd_sc_hd__o31a_1 _15867_ (.A1(_08344_),
    .A2(_08950_),
    .A3(_08954_),
    .B1(_08961_),
    .X(_08962_));
 sky130_fd_sc_hd__xor2_1 _15868_ (.A(_08960_),
    .B(_08962_),
    .X(_08963_));
 sky130_fd_sc_hd__o22a_1 _15869_ (.A1(_08431_),
    .A2(_08344_),
    .B1(_08696_),
    .B2(_08910_),
    .X(_08964_));
 sky130_fd_sc_hd__a21oi_1 _15870_ (.A1(_08912_),
    .A2(_08943_),
    .B1(_08964_),
    .Y(_08965_));
 sky130_fd_sc_hd__nand2_1 _15871_ (.A(_08963_),
    .B(_08965_),
    .Y(_08966_));
 sky130_fd_sc_hd__or2_1 _15872_ (.A(_08963_),
    .B(_08965_),
    .X(_08967_));
 sky130_fd_sc_hd__or2_1 _15873_ (.A(_08956_),
    .B(_08959_),
    .X(_08968_));
 sky130_fd_sc_hd__o2bb2a_1 _15874_ (.A1_N(_08966_),
    .A2_N(_08967_),
    .B1(_08949_),
    .B2(_08968_),
    .X(_08969_));
 sky130_fd_sc_hd__nor3b_1 _15875_ (.A(_08943_),
    .B(_08948_),
    .C_N(_08968_),
    .Y(_08970_));
 sky130_fd_sc_hd__a311o_1 _15876_ (.A1(_08949_),
    .A2(_08956_),
    .A3(_08959_),
    .B1(_08969_),
    .C1(_08970_),
    .X(_08971_));
 sky130_fd_sc_hd__or2_1 _15877_ (.A(_08928_),
    .B(_08929_),
    .X(_08972_));
 sky130_fd_sc_hd__nand2_1 _15878_ (.A(_08930_),
    .B(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__o21a_1 _15879_ (.A1(_08960_),
    .A2(_08962_),
    .B1(_08966_),
    .X(_08974_));
 sky130_fd_sc_hd__xor2_1 _15880_ (.A(_08973_),
    .B(_08974_),
    .X(_08975_));
 sky130_fd_sc_hd__and3_1 _15881_ (.A(_08912_),
    .B(_08943_),
    .C(_08975_),
    .X(_08976_));
 sky130_fd_sc_hd__or2_1 _15882_ (.A(_08932_),
    .B(_08934_),
    .X(_08977_));
 sky130_fd_sc_hd__and2_1 _15883_ (.A(_08935_),
    .B(_08977_),
    .X(_08978_));
 sky130_fd_sc_hd__o21bai_1 _15884_ (.A1(_08973_),
    .A2(_08974_),
    .B1_N(_08976_),
    .Y(_08979_));
 sky130_fd_sc_hd__nor2_1 _15885_ (.A(_08978_),
    .B(_08979_),
    .Y(_08980_));
 sky130_fd_sc_hd__a21oi_1 _15886_ (.A1(_08912_),
    .A2(_08943_),
    .B1(_08975_),
    .Y(_08981_));
 sky130_fd_sc_hd__or3_1 _15887_ (.A(_08976_),
    .B(_08980_),
    .C(_08981_),
    .X(_08982_));
 sky130_fd_sc_hd__a2bb2o_1 _15888_ (.A1_N(_08971_),
    .A2_N(_08982_),
    .B1(_08978_),
    .B2(_08979_),
    .X(_08983_));
 sky130_fd_sc_hd__inv_2 _15889_ (.A(_08898_),
    .Y(_08984_));
 sky130_fd_sc_hd__o22a_1 _15890_ (.A1(_08984_),
    .A2(_08907_),
    .B1(_08938_),
    .B2(_08909_),
    .X(_08985_));
 sky130_fd_sc_hd__xnor2_1 _15891_ (.A(_08916_),
    .B(_08937_),
    .Y(_08986_));
 sky130_fd_sc_hd__a211oi_1 _15892_ (.A1(_08909_),
    .A2(_08938_),
    .B1(_08986_),
    .C1(_08901_),
    .Y(_08987_));
 sky130_fd_sc_hd__and4_1 _15893_ (.A(_08868_),
    .B(_08983_),
    .C(_08985_),
    .D(_08987_),
    .X(_08988_));
 sky130_fd_sc_hd__and2b_1 _15894_ (.A_N(_08906_),
    .B(_08941_),
    .X(_08989_));
 sky130_fd_sc_hd__a21o_1 _15895_ (.A1(_08942_),
    .A2(_08988_),
    .B1(_08989_),
    .X(_08990_));
 sky130_fd_sc_hd__a22o_2 _15896_ (.A1(_08865_),
    .A2(_08903_),
    .B1(_08905_),
    .B2(_08990_),
    .X(_08991_));
 sky130_fd_sc_hd__nor2_1 _15897_ (.A(_08809_),
    .B(_08866_),
    .Y(_08992_));
 sky130_fd_sc_hd__xnor2_2 _15898_ (.A(_08810_),
    .B(_08992_),
    .Y(_08993_));
 sky130_fd_sc_hd__a22o_2 _15899_ (.A1(_08810_),
    .A2(_08866_),
    .B1(_08991_),
    .B2(_08993_),
    .X(_08994_));
 sky130_fd_sc_hd__nand2_1 _15900_ (.A(_08757_),
    .B(_08811_),
    .Y(_08995_));
 sky130_fd_sc_hd__xnor2_2 _15901_ (.A(_08763_),
    .B(_08995_),
    .Y(_08996_));
 sky130_fd_sc_hd__a2bb2o_2 _15902_ (.A1_N(_08763_),
    .A2_N(_08811_),
    .B1(_08994_),
    .B2(_08996_),
    .X(_08997_));
 sky130_fd_sc_hd__nor2_1 _15903_ (.A(_08761_),
    .B(_08764_),
    .Y(_08998_));
 sky130_fd_sc_hd__xnor2_2 _15904_ (.A(_08659_),
    .B(_08998_),
    .Y(_08999_));
 sky130_fd_sc_hd__a22o_2 _15905_ (.A1(_08659_),
    .A2(_08764_),
    .B1(_08997_),
    .B2(_08999_),
    .X(_09000_));
 sky130_fd_sc_hd__a21o_1 _15906_ (.A1(_08555_),
    .A2(_08566_),
    .B1(_08564_),
    .X(_09001_));
 sky130_fd_sc_hd__or2b_1 _15907_ (.A(_08418_),
    .B_N(_08376_),
    .X(_09002_));
 sky130_fd_sc_hd__or3_1 _15908_ (.A(_08150_),
    .B(_08165_),
    .C(_08274_),
    .X(_09003_));
 sky130_fd_sc_hd__or2_1 _15909_ (.A(_08952_),
    .B(_09003_),
    .X(_09004_));
 sky130_fd_sc_hd__clkbuf_4 _15910_ (.A(_08274_),
    .X(_09005_));
 sky130_fd_sc_hd__o22ai_1 _15911_ (.A1(_08151_),
    .A2(_09005_),
    .B1(_08952_),
    .B2(_08166_),
    .Y(_09006_));
 sky130_fd_sc_hd__nand2_1 _15912_ (.A(_09004_),
    .B(_09006_),
    .Y(_09007_));
 sky130_fd_sc_hd__clkbuf_4 _15913_ (.A(_08335_),
    .X(_09008_));
 sky130_fd_sc_hd__nor2_1 _15914_ (.A(_09008_),
    .B(_08553_),
    .Y(_09009_));
 sky130_fd_sc_hd__xnor2_1 _15915_ (.A(_09007_),
    .B(_09009_),
    .Y(_09010_));
 sky130_fd_sc_hd__nor2_1 _15916_ (.A(_08370_),
    .B(_08328_),
    .Y(_09011_));
 sky130_fd_sc_hd__xnor2_1 _15917_ (.A(_08557_),
    .B(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__or2_1 _15918_ (.A(_08253_),
    .B(_08340_),
    .X(_09013_));
 sky130_fd_sc_hd__xnor2_1 _15919_ (.A(_09012_),
    .B(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__nand2_1 _15920_ (.A(_08556_),
    .B(_08557_),
    .Y(_09015_));
 sky130_fd_sc_hd__o31a_1 _15921_ (.A1(_08276_),
    .A2(_08535_),
    .A3(_08558_),
    .B1(_09015_),
    .X(_09016_));
 sky130_fd_sc_hd__nor2_1 _15922_ (.A(_09014_),
    .B(_09016_),
    .Y(_09017_));
 sky130_fd_sc_hd__and2_1 _15923_ (.A(_09014_),
    .B(_09016_),
    .X(_09018_));
 sky130_fd_sc_hd__nor2_1 _15924_ (.A(_09017_),
    .B(_09018_),
    .Y(_09019_));
 sky130_fd_sc_hd__xnor2_1 _15925_ (.A(_09010_),
    .B(_09019_),
    .Y(_09020_));
 sky130_fd_sc_hd__a21o_1 _15926_ (.A1(_08416_),
    .A2(_09002_),
    .B1(_09020_),
    .X(_09021_));
 sky130_fd_sc_hd__nand3_1 _15927_ (.A(_08416_),
    .B(_09002_),
    .C(_09020_),
    .Y(_09022_));
 sky130_fd_sc_hd__nand2_1 _15928_ (.A(_09021_),
    .B(_09022_),
    .Y(_09023_));
 sky130_fd_sc_hd__xnor2_1 _15929_ (.A(_09001_),
    .B(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__a21bo_1 _15930_ (.A1(_08377_),
    .A2(_08385_),
    .B1_N(_08387_),
    .X(_09025_));
 sky130_fd_sc_hd__a21bo_1 _15931_ (.A1(_08432_),
    .A2(_08435_),
    .B1_N(_08430_),
    .X(_09026_));
 sky130_fd_sc_hd__nor2_1 _15932_ (.A(_08516_),
    .B(_08408_),
    .Y(_09027_));
 sky130_fd_sc_hd__o22ai_1 _15933_ (.A1(_08369_),
    .A2(_08408_),
    .B1(_08384_),
    .B2(_08516_),
    .Y(_09028_));
 sky130_fd_sc_hd__a21bo_1 _15934_ (.A1(_08385_),
    .A2(_09027_),
    .B1_N(_09028_),
    .X(_09029_));
 sky130_fd_sc_hd__nor2_1 _15935_ (.A(_08368_),
    .B(_08373_),
    .Y(_09030_));
 sky130_fd_sc_hd__xor2_1 _15936_ (.A(_09029_),
    .B(_09030_),
    .X(_09031_));
 sky130_fd_sc_hd__xnor2_1 _15937_ (.A(_09026_),
    .B(_09031_),
    .Y(_09032_));
 sky130_fd_sc_hd__nand2_1 _15938_ (.A(_09025_),
    .B(_09032_),
    .Y(_09033_));
 sky130_fd_sc_hd__or2_1 _15939_ (.A(_09025_),
    .B(_09032_),
    .X(_09034_));
 sky130_fd_sc_hd__and2_1 _15940_ (.A(_09033_),
    .B(_09034_),
    .X(_09035_));
 sky130_fd_sc_hd__nor2_1 _15941_ (.A(_08910_),
    .B(_08429_),
    .Y(_09036_));
 sky130_fd_sc_hd__clkbuf_4 _15942_ (.A(_08447_),
    .X(_09037_));
 sky130_fd_sc_hd__nor2_1 _15943_ (.A(_08390_),
    .B(_09037_),
    .Y(_09038_));
 sky130_fd_sc_hd__xnor2_2 _15944_ (.A(_09036_),
    .B(_09038_),
    .Y(_09039_));
 sky130_fd_sc_hd__nor2_1 _15945_ (.A(_08434_),
    .B(_08497_),
    .Y(_09040_));
 sky130_fd_sc_hd__xnor2_2 _15946_ (.A(_09039_),
    .B(_09040_),
    .Y(_09041_));
 sky130_fd_sc_hd__nand2_1 _15947_ (.A(\rbzero.wall_tracer.stepDistY[3] ),
    .B(_08338_),
    .Y(_09042_));
 sky130_fd_sc_hd__a21o_1 _15948_ (.A1(_08455_),
    .A2(_09042_),
    .B1(_08357_),
    .X(_09043_));
 sky130_fd_sc_hd__clkbuf_4 _15949_ (.A(_09043_),
    .X(_09044_));
 sky130_fd_sc_hd__buf_6 _15950_ (.A(_08357_),
    .X(_09045_));
 sky130_fd_sc_hd__nand2_8 _15951_ (.A(\rbzero.wall_tracer.stepDistX[3] ),
    .B(_09045_),
    .Y(_09046_));
 sky130_fd_sc_hd__a21oi_2 _15952_ (.A1(_09044_),
    .A2(_09046_),
    .B1(_08441_),
    .Y(_09047_));
 sky130_fd_sc_hd__a21oi_2 _15953_ (.A1(_08462_),
    .A2(_08465_),
    .B1(_08458_),
    .Y(_09048_));
 sky130_fd_sc_hd__or3_1 _15954_ (.A(_08012_),
    .B(_08015_),
    .C(_08450_),
    .X(_09049_));
 sky130_fd_sc_hd__o21ai_1 _15955_ (.A1(_08012_),
    .A2(_08450_),
    .B1(_08015_),
    .Y(_09050_));
 sky130_fd_sc_hd__a31o_1 _15956_ (.A1(_08148_),
    .A2(_09049_),
    .A3(_09050_),
    .B1(_08454_),
    .X(_09051_));
 sky130_fd_sc_hd__nand2_1 _15957_ (.A(\rbzero.wall_tracer.stepDistY[5] ),
    .B(_08338_),
    .Y(_09052_));
 sky130_fd_sc_hd__a21o_2 _15958_ (.A1(_09051_),
    .A2(_09052_),
    .B1(_08357_),
    .X(_09053_));
 sky130_fd_sc_hd__nor2_1 _15959_ (.A(_08461_),
    .B(_09053_),
    .Y(_09054_));
 sky130_fd_sc_hd__xor2_2 _15960_ (.A(_09048_),
    .B(_09054_),
    .X(_09055_));
 sky130_fd_sc_hd__xor2_2 _15961_ (.A(_09047_),
    .B(_09055_),
    .X(_09056_));
 sky130_fd_sc_hd__or3_1 _15962_ (.A(_09043_),
    .B(_08581_),
    .C(_08467_),
    .X(_09057_));
 sky130_fd_sc_hd__a21bo_1 _15963_ (.A1(_08448_),
    .A2(_08468_),
    .B1_N(_09057_),
    .X(_09058_));
 sky130_fd_sc_hd__xor2_2 _15964_ (.A(_09056_),
    .B(_09058_),
    .X(_09059_));
 sky130_fd_sc_hd__xnor2_2 _15965_ (.A(_09041_),
    .B(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__nor2_1 _15966_ (.A(_08469_),
    .B(_08478_),
    .Y(_09061_));
 sky130_fd_sc_hd__a21o_1 _15967_ (.A1(_08436_),
    .A2(_08479_),
    .B1(_09061_),
    .X(_09062_));
 sky130_fd_sc_hd__xnor2_2 _15968_ (.A(_09060_),
    .B(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__xnor2_2 _15969_ (.A(_09035_),
    .B(_09063_),
    .Y(_09064_));
 sky130_fd_sc_hd__or2b_1 _15970_ (.A(_08480_),
    .B_N(_08493_),
    .X(_09065_));
 sky130_fd_sc_hd__a21boi_1 _15971_ (.A1(_08419_),
    .A2(_08494_),
    .B1_N(_09065_),
    .Y(_09066_));
 sky130_fd_sc_hd__xor2_1 _15972_ (.A(_09064_),
    .B(_09066_),
    .X(_09067_));
 sky130_fd_sc_hd__xnor2_1 _15973_ (.A(_09024_),
    .B(_09067_),
    .Y(_09068_));
 sky130_fd_sc_hd__and2b_1 _15974_ (.A_N(_08495_),
    .B(_08527_),
    .X(_09069_));
 sky130_fd_sc_hd__a21oi_1 _15975_ (.A1(_08528_),
    .A2(_08571_),
    .B1(_09069_),
    .Y(_09070_));
 sky130_fd_sc_hd__nor2_1 _15976_ (.A(_09068_),
    .B(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__nand2_1 _15977_ (.A(_09068_),
    .B(_09070_),
    .Y(_09072_));
 sky130_fd_sc_hd__and2b_1 _15978_ (.A_N(_09071_),
    .B(_09072_),
    .X(_09073_));
 sky130_fd_sc_hd__or2b_1 _15979_ (.A(_08570_),
    .B_N(_08546_),
    .X(_09074_));
 sky130_fd_sc_hd__a21bo_1 _15980_ (.A1(_08549_),
    .A2(_08550_),
    .B1_N(_08552_),
    .X(_09075_));
 sky130_fd_sc_hd__nand2_4 _15981_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08149_),
    .Y(_09076_));
 sky130_fd_sc_hd__or2_1 _15982_ (.A(_08164_),
    .B(_09076_),
    .X(_09077_));
 sky130_fd_sc_hd__nor2_1 _15983_ (.A(_08619_),
    .B(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__clkbuf_4 _15984_ (.A(_09076_),
    .X(_09079_));
 sky130_fd_sc_hd__o22a_1 _15985_ (.A1(_08304_),
    .A2(_08618_),
    .B1(_09079_),
    .B2(_08616_),
    .X(_09080_));
 sky130_fd_sc_hd__or2_1 _15986_ (.A(_09078_),
    .B(_09080_),
    .X(_09081_));
 sky130_fd_sc_hd__xnor2_1 _15987_ (.A(_09075_),
    .B(_09081_),
    .Y(_09082_));
 sky130_fd_sc_hd__nand2_1 _15988_ (.A(_08622_),
    .B(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__or2_1 _15989_ (.A(_08622_),
    .B(_09082_),
    .X(_09084_));
 sky130_fd_sc_hd__nand2_1 _15990_ (.A(_09083_),
    .B(_09084_),
    .Y(_09085_));
 sky130_fd_sc_hd__a21oi_4 _15991_ (.A1(_08568_),
    .A2(_09074_),
    .B1(_09085_),
    .Y(_09086_));
 sky130_fd_sc_hd__and3_1 _15992_ (.A(_08568_),
    .B(_09074_),
    .C(_09085_),
    .X(_09087_));
 sky130_fd_sc_hd__nor2_1 _15993_ (.A(_09086_),
    .B(_09087_),
    .Y(_09088_));
 sky130_fd_sc_hd__xnor2_2 _15994_ (.A(_09073_),
    .B(_09088_),
    .Y(_09089_));
 sky130_fd_sc_hd__nor2_1 _15995_ (.A(_08572_),
    .B(_08613_),
    .Y(_09090_));
 sky130_fd_sc_hd__a21oi_2 _15996_ (.A1(_08614_),
    .A2(_08627_),
    .B1(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__xor2_2 _15997_ (.A(_09089_),
    .B(_09091_),
    .X(_09092_));
 sky130_fd_sc_hd__xnor2_1 _15998_ (.A(_08625_),
    .B(_09092_),
    .Y(_09093_));
 sky130_fd_sc_hd__or2b_1 _15999_ (.A(_08367_),
    .B_N(_08658_),
    .X(_09094_));
 sky130_fd_sc_hd__o21a_1 _16000_ (.A1(_08628_),
    .A2(_08657_),
    .B1(_09094_),
    .X(_09095_));
 sky130_fd_sc_hd__xor2_1 _16001_ (.A(_09093_),
    .B(_09095_),
    .X(_09096_));
 sky130_fd_sc_hd__and2_1 _16002_ (.A(_08659_),
    .B(_08761_),
    .X(_09097_));
 sky130_fd_sc_hd__nand2_1 _16003_ (.A(_09096_),
    .B(_09097_),
    .Y(_09098_));
 sky130_fd_sc_hd__or2_1 _16004_ (.A(_09096_),
    .B(_09097_),
    .X(_09099_));
 sky130_fd_sc_hd__and2_2 _16005_ (.A(_09098_),
    .B(_09099_),
    .X(_09100_));
 sky130_fd_sc_hd__xor2_4 _16006_ (.A(_09000_),
    .B(_09100_),
    .X(_09101_));
 sky130_fd_sc_hd__clkinv_2 _16007_ (.A(\rbzero.debug_overlay.playerX[-6] ),
    .Y(_09102_));
 sky130_fd_sc_hd__mux2_1 _16008_ (.A0(_08220_),
    .A1(_09102_),
    .S(_08138_),
    .X(_09103_));
 sky130_fd_sc_hd__xnor2_1 _16009_ (.A(_09101_),
    .B(_09103_),
    .Y(_09104_));
 sky130_fd_sc_hd__xor2_4 _16010_ (.A(_08997_),
    .B(_08999_),
    .X(_09105_));
 sky130_fd_sc_hd__mux2_1 _16011_ (.A0(\rbzero.debug_overlay.playerY[-7] ),
    .A1(\rbzero.debug_overlay.playerX[-7] ),
    .S(_08138_),
    .X(_09106_));
 sky130_fd_sc_hd__or2_1 _16012_ (.A(_09105_),
    .B(_09106_),
    .X(_09107_));
 sky130_fd_sc_hd__xor2_4 _16013_ (.A(_08991_),
    .B(_08993_),
    .X(_09108_));
 sky130_fd_sc_hd__mux2_1 _16014_ (.A0(\rbzero.debug_overlay.playerY[-9] ),
    .A1(\rbzero.debug_overlay.playerX[-9] ),
    .S(_08138_),
    .X(_09109_));
 sky130_fd_sc_hd__mux2_1 _16015_ (.A0(\rbzero.debug_overlay.playerY[-8] ),
    .A1(\rbzero.debug_overlay.playerX[-8] ),
    .S(_04464_),
    .X(_09110_));
 sky130_fd_sc_hd__xor2_4 _16016_ (.A(_08994_),
    .B(_08996_),
    .X(_09111_));
 sky130_fd_sc_hd__or2_1 _16017_ (.A(_09110_),
    .B(_09111_),
    .X(_09112_));
 sky130_fd_sc_hd__and2_1 _16018_ (.A(_09110_),
    .B(_09111_),
    .X(_09113_));
 sky130_fd_sc_hd__a31o_1 _16019_ (.A1(_09108_),
    .A2(_09109_),
    .A3(_09112_),
    .B1(_09113_),
    .X(_09114_));
 sky130_fd_sc_hd__and2_1 _16020_ (.A(_09105_),
    .B(_09106_),
    .X(_09115_));
 sky130_fd_sc_hd__a21o_1 _16021_ (.A1(_09107_),
    .A2(_09114_),
    .B1(_09115_),
    .X(_09116_));
 sky130_fd_sc_hd__xnor2_1 _16022_ (.A(_09104_),
    .B(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__clkbuf_4 _16023_ (.A(_08218_),
    .X(_09118_));
 sky130_fd_sc_hd__buf_2 _16024_ (.A(_09118_),
    .X(_09119_));
 sky130_fd_sc_hd__mux2_1 _16025_ (.A0(_06087_),
    .A1(_09119_),
    .S(_08395_),
    .X(_09120_));
 sky130_fd_sc_hd__buf_2 _16026_ (.A(_09120_),
    .X(_09121_));
 sky130_fd_sc_hd__and2_1 _16027_ (.A(_09117_),
    .B(_09121_),
    .X(_09122_));
 sky130_fd_sc_hd__nor2_1 _16028_ (.A(_09117_),
    .B(_09121_),
    .Y(_09123_));
 sky130_fd_sc_hd__or3_2 _16029_ (.A(_08148_),
    .B(_09122_),
    .C(_09123_),
    .X(_09124_));
 sky130_fd_sc_hd__o211a_1 _16030_ (.A1(\rbzero.texu_hot[0] ),
    .A2(_08145_),
    .B1(_09124_),
    .C1(_08085_),
    .X(_00466_));
 sky130_fd_sc_hd__a21boi_2 _16031_ (.A1(_09000_),
    .A2(_09100_),
    .B1_N(_09098_),
    .Y(_09125_));
 sky130_fd_sc_hd__or2_2 _16032_ (.A(_09093_),
    .B(_09095_),
    .X(_09126_));
 sky130_fd_sc_hd__or2b_1 _16033_ (.A(_09023_),
    .B_N(_09001_),
    .X(_09127_));
 sky130_fd_sc_hd__or3_1 _16034_ (.A(_09008_),
    .B(_08553_),
    .C(_09007_),
    .X(_09128_));
 sky130_fd_sc_hd__nor2_1 _16035_ (.A(_08335_),
    .B(_08618_),
    .Y(_09129_));
 sky130_fd_sc_hd__xnor2_1 _16036_ (.A(_09077_),
    .B(_09129_),
    .Y(_09130_));
 sky130_fd_sc_hd__nand2_4 _16037_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08475_),
    .Y(_09131_));
 sky130_fd_sc_hd__nor2_1 _16038_ (.A(_08171_),
    .B(_09131_),
    .Y(_09132_));
 sky130_fd_sc_hd__xnor2_1 _16039_ (.A(_09130_),
    .B(_09132_),
    .Y(_09133_));
 sky130_fd_sc_hd__nand3_1 _16040_ (.A(_09004_),
    .B(_09128_),
    .C(_09133_),
    .Y(_09134_));
 sky130_fd_sc_hd__a21o_1 _16041_ (.A1(_09004_),
    .A2(_09128_),
    .B1(_09133_),
    .X(_09135_));
 sky130_fd_sc_hd__nand2_1 _16042_ (.A(_09134_),
    .B(_09135_),
    .Y(_09136_));
 sky130_fd_sc_hd__and2b_1 _16043_ (.A_N(_09081_),
    .B(_09075_),
    .X(_09137_));
 sky130_fd_sc_hd__nor2_1 _16044_ (.A(_09078_),
    .B(_09137_),
    .Y(_09138_));
 sky130_fd_sc_hd__xnor2_1 _16045_ (.A(_09136_),
    .B(_09138_),
    .Y(_09139_));
 sky130_fd_sc_hd__a21oi_1 _16046_ (.A1(_09021_),
    .A2(_09127_),
    .B1(_09139_),
    .Y(_09140_));
 sky130_fd_sc_hd__and3_1 _16047_ (.A(_09021_),
    .B(_09127_),
    .C(_09139_),
    .X(_09141_));
 sky130_fd_sc_hd__nor2_1 _16048_ (.A(_09140_),
    .B(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__xnor2_1 _16049_ (.A(_09083_),
    .B(_09142_),
    .Y(_09143_));
 sky130_fd_sc_hd__a21o_1 _16050_ (.A1(_09010_),
    .A2(_09019_),
    .B1(_09017_),
    .X(_09144_));
 sky130_fd_sc_hd__or2b_1 _16051_ (.A(_09031_),
    .B_N(_09026_),
    .X(_09145_));
 sky130_fd_sc_hd__clkbuf_4 _16052_ (.A(_08847_),
    .X(_09146_));
 sky130_fd_sc_hd__o22ai_1 _16053_ (.A1(_08152_),
    .A2(_08847_),
    .B1(_09005_),
    .B2(_08166_),
    .Y(_09147_));
 sky130_fd_sc_hd__o21ai_1 _16054_ (.A1(_09146_),
    .A2(_09003_),
    .B1(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__nor2_1 _16055_ (.A(_08952_),
    .B(_08553_),
    .Y(_09149_));
 sky130_fd_sc_hd__xnor2_1 _16056_ (.A(_09148_),
    .B(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__or2_1 _16057_ (.A(_08370_),
    .B(_08325_),
    .X(_09151_));
 sky130_fd_sc_hd__nor2_1 _16058_ (.A(_08368_),
    .B(_08328_),
    .Y(_09152_));
 sky130_fd_sc_hd__xnor2_1 _16059_ (.A(_09151_),
    .B(_09152_),
    .Y(_09153_));
 sky130_fd_sc_hd__nor2_1 _16060_ (.A(_08235_),
    .B(_08340_),
    .Y(_09154_));
 sky130_fd_sc_hd__xnor2_1 _16061_ (.A(_09153_),
    .B(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__nand2_1 _16062_ (.A(_08557_),
    .B(_09011_),
    .Y(_09156_));
 sky130_fd_sc_hd__o31a_1 _16063_ (.A1(_08253_),
    .A2(_08535_),
    .A3(_09012_),
    .B1(_09156_),
    .X(_09157_));
 sky130_fd_sc_hd__nor2_1 _16064_ (.A(_09155_),
    .B(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__and2_1 _16065_ (.A(_09155_),
    .B(_09157_),
    .X(_09159_));
 sky130_fd_sc_hd__nor2_1 _16066_ (.A(_09158_),
    .B(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__xnor2_1 _16067_ (.A(_09150_),
    .B(_09160_),
    .Y(_09161_));
 sky130_fd_sc_hd__a21o_1 _16068_ (.A1(_09145_),
    .A2(_09033_),
    .B1(_09161_),
    .X(_09162_));
 sky130_fd_sc_hd__nand3_1 _16069_ (.A(_09145_),
    .B(_09033_),
    .C(_09161_),
    .Y(_09163_));
 sky130_fd_sc_hd__nand2_1 _16070_ (.A(_09162_),
    .B(_09163_),
    .Y(_09164_));
 sky130_fd_sc_hd__xnor2_1 _16071_ (.A(_09144_),
    .B(_09164_),
    .Y(_09165_));
 sky130_fd_sc_hd__a22o_1 _16072_ (.A1(_08385_),
    .A2(_09027_),
    .B1(_09028_),
    .B2(_09030_),
    .X(_09166_));
 sky130_fd_sc_hd__clkbuf_4 _16073_ (.A(_08434_),
    .X(_09167_));
 sky130_fd_sc_hd__nand2_1 _16074_ (.A(_09036_),
    .B(_09038_),
    .Y(_09168_));
 sky130_fd_sc_hd__o31a_1 _16075_ (.A1(_09167_),
    .A2(_08497_),
    .A3(_09039_),
    .B1(_09168_),
    .X(_09169_));
 sky130_fd_sc_hd__nor2_2 _16076_ (.A(_08369_),
    .B(_08497_),
    .Y(_09170_));
 sky130_fd_sc_hd__xor2_1 _16077_ (.A(_09027_),
    .B(_09170_),
    .X(_09171_));
 sky130_fd_sc_hd__nor2_1 _16078_ (.A(_08373_),
    .B(_08384_),
    .Y(_09172_));
 sky130_fd_sc_hd__xnor2_1 _16079_ (.A(_09171_),
    .B(_09172_),
    .Y(_09173_));
 sky130_fd_sc_hd__xnor2_1 _16080_ (.A(_09169_),
    .B(_09173_),
    .Y(_09174_));
 sky130_fd_sc_hd__xnor2_2 _16081_ (.A(_09166_),
    .B(_09174_),
    .Y(_09175_));
 sky130_fd_sc_hd__buf_2 _16082_ (.A(_08429_),
    .X(_09176_));
 sky130_fd_sc_hd__nor2_1 _16083_ (.A(_08434_),
    .B(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__or2_1 _16084_ (.A(_08410_),
    .B(_08447_),
    .X(_09178_));
 sky130_fd_sc_hd__a21oi_1 _16085_ (.A1(_09044_),
    .A2(_09046_),
    .B1(_08390_),
    .Y(_09179_));
 sky130_fd_sc_hd__xnor2_1 _16086_ (.A(_09178_),
    .B(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__and2_1 _16087_ (.A(_09177_),
    .B(_09180_),
    .X(_09181_));
 sky130_fd_sc_hd__nor2_1 _16088_ (.A(_09177_),
    .B(_09180_),
    .Y(_09182_));
 sky130_fd_sc_hd__nor2_1 _16089_ (.A(_09181_),
    .B(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__nand2_4 _16090_ (.A(\rbzero.wall_tracer.stepDistX[4] ),
    .B(_08357_),
    .Y(_09184_));
 sky130_fd_sc_hd__and2_1 _16091_ (.A(_08466_),
    .B(_09184_),
    .X(_09185_));
 sky130_fd_sc_hd__buf_2 _16092_ (.A(_09185_),
    .X(_09186_));
 sky130_fd_sc_hd__o31a_1 _16093_ (.A1(_08012_),
    .A2(_08015_),
    .A3(_08450_),
    .B1(_08018_),
    .X(_09187_));
 sky130_fd_sc_hd__or2_1 _16094_ (.A(_08015_),
    .B(_08018_),
    .X(_09188_));
 sky130_fd_sc_hd__nor3_1 _16095_ (.A(_08012_),
    .B(_08450_),
    .C(_09188_),
    .Y(_09189_));
 sky130_fd_sc_hd__a31oi_4 _16096_ (.A1(_08144_),
    .A2(_08452_),
    .A3(_08453_),
    .B1(_08405_),
    .Y(_09190_));
 sky130_fd_sc_hd__o31ai_4 _16097_ (.A1(_08145_),
    .A2(_09187_),
    .A3(_09189_),
    .B1(_09190_),
    .Y(_09191_));
 sky130_fd_sc_hd__or3_2 _16098_ (.A(_08042_),
    .B(_08338_),
    .C(_09191_),
    .X(_09192_));
 sky130_fd_sc_hd__nor3_1 _16099_ (.A(_08461_),
    .B(_09053_),
    .C(_09192_),
    .Y(_09193_));
 sky130_fd_sc_hd__nand2_1 _16100_ (.A(\rbzero.wall_tracer.stepDistY[6] ),
    .B(_08405_),
    .Y(_09194_));
 sky130_fd_sc_hd__a21o_4 _16101_ (.A1(_09194_),
    .A2(_09191_),
    .B1(_09045_),
    .X(_09195_));
 sky130_fd_sc_hd__o22a_1 _16102_ (.A1(_08581_),
    .A2(_09053_),
    .B1(_09195_),
    .B2(_08461_),
    .X(_09196_));
 sky130_fd_sc_hd__or4_1 _16103_ (.A(_08441_),
    .B(_09186_),
    .C(_09193_),
    .D(_09196_),
    .X(_09197_));
 sky130_fd_sc_hd__o22ai_1 _16104_ (.A1(_08950_),
    .A2(_09186_),
    .B1(_09193_),
    .B2(_09196_),
    .Y(_09198_));
 sky130_fd_sc_hd__nand2_1 _16105_ (.A(_09197_),
    .B(_09198_),
    .Y(_09199_));
 sky130_fd_sc_hd__nand2_1 _16106_ (.A(_09048_),
    .B(_09054_),
    .Y(_09200_));
 sky130_fd_sc_hd__a21bo_1 _16107_ (.A1(_09047_),
    .A2(_09055_),
    .B1_N(_09200_),
    .X(_09201_));
 sky130_fd_sc_hd__xnor2_2 _16108_ (.A(_09199_),
    .B(_09201_),
    .Y(_09202_));
 sky130_fd_sc_hd__xnor2_2 _16109_ (.A(_09183_),
    .B(_09202_),
    .Y(_09203_));
 sky130_fd_sc_hd__nand2_1 _16110_ (.A(_09056_),
    .B(_09058_),
    .Y(_09204_));
 sky130_fd_sc_hd__a21bo_1 _16111_ (.A1(_09041_),
    .A2(_09059_),
    .B1_N(_09204_),
    .X(_09205_));
 sky130_fd_sc_hd__xnor2_2 _16112_ (.A(_09203_),
    .B(_09205_),
    .Y(_09206_));
 sky130_fd_sc_hd__xnor2_2 _16113_ (.A(_09175_),
    .B(_09206_),
    .Y(_09207_));
 sky130_fd_sc_hd__and2b_1 _16114_ (.A_N(_09060_),
    .B(_09062_),
    .X(_09208_));
 sky130_fd_sc_hd__a21oi_1 _16115_ (.A1(_09035_),
    .A2(_09063_),
    .B1(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__xor2_1 _16116_ (.A(_09207_),
    .B(_09209_),
    .X(_09210_));
 sky130_fd_sc_hd__xnor2_1 _16117_ (.A(_09165_),
    .B(_09210_),
    .Y(_09211_));
 sky130_fd_sc_hd__nor2_1 _16118_ (.A(_09064_),
    .B(_09066_),
    .Y(_09212_));
 sky130_fd_sc_hd__a21oi_1 _16119_ (.A1(_09024_),
    .A2(_09067_),
    .B1(_09212_),
    .Y(_09213_));
 sky130_fd_sc_hd__nor2_1 _16120_ (.A(_09211_),
    .B(_09213_),
    .Y(_09214_));
 sky130_fd_sc_hd__and2_1 _16121_ (.A(_09211_),
    .B(_09213_),
    .X(_09215_));
 sky130_fd_sc_hd__nor2_1 _16122_ (.A(_09214_),
    .B(_09215_),
    .Y(_09216_));
 sky130_fd_sc_hd__xnor2_1 _16123_ (.A(_09143_),
    .B(_09216_),
    .Y(_09217_));
 sky130_fd_sc_hd__a21oi_1 _16124_ (.A1(_09072_),
    .A2(_09088_),
    .B1(_09071_),
    .Y(_09218_));
 sky130_fd_sc_hd__nor2_1 _16125_ (.A(_09217_),
    .B(_09218_),
    .Y(_09219_));
 sky130_fd_sc_hd__nand2_1 _16126_ (.A(_09217_),
    .B(_09218_),
    .Y(_09220_));
 sky130_fd_sc_hd__and2b_1 _16127_ (.A_N(_09219_),
    .B(_09220_),
    .X(_09221_));
 sky130_fd_sc_hd__xnor2_4 _16128_ (.A(_09086_),
    .B(_09221_),
    .Y(_09222_));
 sky130_fd_sc_hd__nor2_1 _16129_ (.A(_09089_),
    .B(_09091_),
    .Y(_09223_));
 sky130_fd_sc_hd__a21oi_4 _16130_ (.A1(_08625_),
    .A2(_09092_),
    .B1(_09223_),
    .Y(_09224_));
 sky130_fd_sc_hd__xnor2_4 _16131_ (.A(_09222_),
    .B(_09224_),
    .Y(_09225_));
 sky130_fd_sc_hd__xor2_4 _16132_ (.A(_09126_),
    .B(_09225_),
    .X(_09226_));
 sky130_fd_sc_hd__xnor2_4 _16133_ (.A(_09125_),
    .B(_09226_),
    .Y(_09227_));
 sky130_fd_sc_hd__mux2_1 _16134_ (.A0(\rbzero.debug_overlay.playerY[-5] ),
    .A1(\rbzero.debug_overlay.playerX[-5] ),
    .S(_08138_),
    .X(_09228_));
 sky130_fd_sc_hd__xnor2_1 _16135_ (.A(_09227_),
    .B(_09228_),
    .Y(_09229_));
 sky130_fd_sc_hd__and2b_1 _16136_ (.A_N(_09103_),
    .B(_09101_),
    .X(_09230_));
 sky130_fd_sc_hd__a21oi_1 _16137_ (.A1(_09104_),
    .A2(_09116_),
    .B1(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__or2_1 _16138_ (.A(_09229_),
    .B(_09231_),
    .X(_09232_));
 sky130_fd_sc_hd__nand2_1 _16139_ (.A(_09229_),
    .B(_09231_),
    .Y(_09233_));
 sky130_fd_sc_hd__nand2_1 _16140_ (.A(_09232_),
    .B(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__and2_1 _16141_ (.A(_09121_),
    .B(_09234_),
    .X(_09235_));
 sky130_fd_sc_hd__nor2_1 _16142_ (.A(_09121_),
    .B(_09234_),
    .Y(_09236_));
 sky130_fd_sc_hd__or3_2 _16143_ (.A(_08148_),
    .B(_09235_),
    .C(_09236_),
    .X(_09237_));
 sky130_fd_sc_hd__o211a_1 _16144_ (.A1(\rbzero.texu_hot[1] ),
    .A2(_08145_),
    .B1(_09237_),
    .C1(_08085_),
    .X(_00467_));
 sky130_fd_sc_hd__nand2_1 _16145_ (.A(_09227_),
    .B(_09228_),
    .Y(_09238_));
 sky130_fd_sc_hd__a31o_1 _16146_ (.A1(_08622_),
    .A2(_09082_),
    .A3(_09142_),
    .B1(_09140_),
    .X(_09239_));
 sky130_fd_sc_hd__or2b_1 _16147_ (.A(_09164_),
    .B_N(_09144_),
    .X(_09240_));
 sky130_fd_sc_hd__nand2_1 _16148_ (.A(_09162_),
    .B(_09240_),
    .Y(_09241_));
 sky130_fd_sc_hd__nand2_4 _16149_ (.A(\rbzero.wall_tracer.visualWallDist[7] ),
    .B(_08475_),
    .Y(_09242_));
 sky130_fd_sc_hd__buf_4 _16150_ (.A(_09242_),
    .X(_09243_));
 sky130_fd_sc_hd__nor2_2 _16151_ (.A(_08616_),
    .B(_09243_),
    .Y(_09244_));
 sky130_fd_sc_hd__or3_1 _16152_ (.A(_09008_),
    .B(_08618_),
    .C(_09077_),
    .X(_09245_));
 sky130_fd_sc_hd__a21bo_1 _16153_ (.A1(_09130_),
    .A2(_09132_),
    .B1_N(_09245_),
    .X(_09246_));
 sky130_fd_sc_hd__inv_2 _16154_ (.A(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__nor2_1 _16155_ (.A(_08335_),
    .B(_09076_),
    .Y(_09248_));
 sky130_fd_sc_hd__nor2_1 _16156_ (.A(_08296_),
    .B(_08617_),
    .Y(_09249_));
 sky130_fd_sc_hd__xnor2_1 _16157_ (.A(_09248_),
    .B(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__or3_1 _16158_ (.A(_08304_),
    .B(_09131_),
    .C(_09250_),
    .X(_09251_));
 sky130_fd_sc_hd__buf_4 _16159_ (.A(_09131_),
    .X(_09252_));
 sky130_fd_sc_hd__o21ai_1 _16160_ (.A1(_08304_),
    .A2(_09252_),
    .B1(_09250_),
    .Y(_09253_));
 sky130_fd_sc_hd__nand2_1 _16161_ (.A(_09251_),
    .B(_09253_),
    .Y(_09254_));
 sky130_fd_sc_hd__nor2_1 _16162_ (.A(_09146_),
    .B(_09003_),
    .Y(_09255_));
 sky130_fd_sc_hd__a21o_1 _16163_ (.A1(_09147_),
    .A2(_09149_),
    .B1(_09255_),
    .X(_09256_));
 sky130_fd_sc_hd__or2b_1 _16164_ (.A(_09254_),
    .B_N(_09256_),
    .X(_09257_));
 sky130_fd_sc_hd__or2b_1 _16165_ (.A(_09256_),
    .B_N(_09254_),
    .X(_09258_));
 sky130_fd_sc_hd__nand2_1 _16166_ (.A(_09257_),
    .B(_09258_),
    .Y(_09259_));
 sky130_fd_sc_hd__xnor2_1 _16167_ (.A(_09247_),
    .B(_09259_),
    .Y(_09260_));
 sky130_fd_sc_hd__inv_2 _16168_ (.A(_09135_),
    .Y(_09261_));
 sky130_fd_sc_hd__o21ai_1 _16169_ (.A1(_09078_),
    .A2(_09261_),
    .B1(_09134_),
    .Y(_09262_));
 sky130_fd_sc_hd__xor2_1 _16170_ (.A(_09260_),
    .B(_09262_),
    .X(_09263_));
 sky130_fd_sc_hd__xnor2_1 _16171_ (.A(_09244_),
    .B(_09263_),
    .Y(_09264_));
 sky130_fd_sc_hd__xor2_1 _16172_ (.A(_09241_),
    .B(_09264_),
    .X(_09265_));
 sky130_fd_sc_hd__or3b_1 _16173_ (.A(_09081_),
    .B(_09136_),
    .C_N(_09075_),
    .X(_09266_));
 sky130_fd_sc_hd__xor2_1 _16174_ (.A(_09265_),
    .B(_09266_),
    .X(_09267_));
 sky130_fd_sc_hd__a21o_1 _16175_ (.A1(_09150_),
    .A2(_09160_),
    .B1(_09158_),
    .X(_09268_));
 sky130_fd_sc_hd__or2b_1 _16176_ (.A(_09174_),
    .B_N(_09166_),
    .X(_09269_));
 sky130_fd_sc_hd__o21ai_1 _16177_ (.A1(_09169_),
    .A2(_09173_),
    .B1(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__or4_1 _16178_ (.A(_08151_),
    .B(_08165_),
    .C(_08731_),
    .D(_08847_),
    .X(_09271_));
 sky130_fd_sc_hd__o22ai_1 _16179_ (.A1(_08151_),
    .A2(_08731_),
    .B1(_08847_),
    .B2(_08166_),
    .Y(_09272_));
 sky130_fd_sc_hd__nand2_1 _16180_ (.A(_09271_),
    .B(_09272_),
    .Y(_09273_));
 sky130_fd_sc_hd__nor2_1 _16181_ (.A(_09005_),
    .B(_08553_),
    .Y(_09274_));
 sky130_fd_sc_hd__xnor2_1 _16182_ (.A(_09273_),
    .B(_09274_),
    .Y(_09275_));
 sky130_fd_sc_hd__nor2_1 _16183_ (.A(_08327_),
    .B(_08384_),
    .Y(_09276_));
 sky130_fd_sc_hd__o22a_1 _16184_ (.A1(_08368_),
    .A2(_08327_),
    .B1(_08384_),
    .B2(_08813_),
    .X(_09277_));
 sky130_fd_sc_hd__a21o_1 _16185_ (.A1(_09152_),
    .A2(_09276_),
    .B1(_09277_),
    .X(_09278_));
 sky130_fd_sc_hd__or2_1 _16186_ (.A(_08370_),
    .B(_08340_),
    .X(_09279_));
 sky130_fd_sc_hd__xnor2_1 _16187_ (.A(_09278_),
    .B(_09279_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand2_1 _16188_ (.A(_09153_),
    .B(_09154_),
    .Y(_09281_));
 sky130_fd_sc_hd__o31a_1 _16189_ (.A1(_08368_),
    .A2(_08814_),
    .A3(_09151_),
    .B1(_09281_),
    .X(_09282_));
 sky130_fd_sc_hd__xor2_1 _16190_ (.A(_09280_),
    .B(_09282_),
    .X(_09283_));
 sky130_fd_sc_hd__nand2_1 _16191_ (.A(_09275_),
    .B(_09283_),
    .Y(_09284_));
 sky130_fd_sc_hd__or2_1 _16192_ (.A(_09275_),
    .B(_09283_),
    .X(_09285_));
 sky130_fd_sc_hd__and2_1 _16193_ (.A(_09284_),
    .B(_09285_),
    .X(_09286_));
 sky130_fd_sc_hd__xnor2_1 _16194_ (.A(_09270_),
    .B(_09286_),
    .Y(_09287_));
 sky130_fd_sc_hd__xnor2_1 _16195_ (.A(_09268_),
    .B(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__a22o_1 _16196_ (.A1(_09027_),
    .A2(_09170_),
    .B1(_09171_),
    .B2(_09172_),
    .X(_09289_));
 sky130_fd_sc_hd__a21oi_2 _16197_ (.A1(_09043_),
    .A2(_09046_),
    .B1(_08910_),
    .Y(_09290_));
 sky130_fd_sc_hd__nand2_1 _16198_ (.A(_09038_),
    .B(_09290_),
    .Y(_09291_));
 sky130_fd_sc_hd__inv_2 _16199_ (.A(_09291_),
    .Y(_09292_));
 sky130_fd_sc_hd__nor2_1 _16200_ (.A(_08516_),
    .B(_08429_),
    .Y(_09293_));
 sky130_fd_sc_hd__o22a_1 _16201_ (.A1(_08516_),
    .A2(_08400_),
    .B1(_08429_),
    .B2(_08369_),
    .X(_09294_));
 sky130_fd_sc_hd__a21o_1 _16202_ (.A1(_09170_),
    .A2(_09293_),
    .B1(_09294_),
    .X(_09295_));
 sky130_fd_sc_hd__nor2_1 _16203_ (.A(_08373_),
    .B(_08409_),
    .Y(_09296_));
 sky130_fd_sc_hd__xnor2_1 _16204_ (.A(_09295_),
    .B(_09296_),
    .Y(_09297_));
 sky130_fd_sc_hd__o21ai_1 _16205_ (.A1(_09292_),
    .A2(_09181_),
    .B1(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__a211o_1 _16206_ (.A1(_09177_),
    .A2(_09180_),
    .B1(_09297_),
    .C1(_09292_),
    .X(_09299_));
 sky130_fd_sc_hd__and2_1 _16207_ (.A(_09298_),
    .B(_09299_),
    .X(_09300_));
 sky130_fd_sc_hd__xor2_1 _16208_ (.A(_09289_),
    .B(_09300_),
    .X(_09301_));
 sky130_fd_sc_hd__nor2_1 _16209_ (.A(_08434_),
    .B(_09037_),
    .Y(_09302_));
 sky130_fd_sc_hd__a21oi_2 _16210_ (.A1(_08466_),
    .A2(_09184_),
    .B1(_08390_),
    .Y(_09303_));
 sky130_fd_sc_hd__xor2_2 _16211_ (.A(_09290_),
    .B(_09303_),
    .X(_09304_));
 sky130_fd_sc_hd__xor2_2 _16212_ (.A(_09302_),
    .B(_09304_),
    .X(_09305_));
 sky130_fd_sc_hd__nand2_4 _16213_ (.A(\rbzero.wall_tracer.stepDistX[5] ),
    .B(_09045_),
    .Y(_09306_));
 sky130_fd_sc_hd__a21oi_2 _16214_ (.A1(_09053_),
    .A2(_09306_),
    .B1(_08441_),
    .Y(_09307_));
 sky130_fd_sc_hd__nor4_1 _16215_ (.A(_08012_),
    .B(_08023_),
    .C(_08450_),
    .D(_09188_),
    .Y(_09308_));
 sky130_fd_sc_hd__o31a_1 _16216_ (.A1(_08012_),
    .A2(_08450_),
    .A3(_09188_),
    .B1(_08023_),
    .X(_09309_));
 sky130_fd_sc_hd__o31a_2 _16217_ (.A1(_08145_),
    .A2(_09308_),
    .A3(_09309_),
    .B1(_09190_),
    .X(_09310_));
 sky130_fd_sc_hd__and3_1 _16218_ (.A(\rbzero.wall_tracer.visualWallDist[-11] ),
    .B(_08149_),
    .C(_09310_),
    .X(_09311_));
 sky130_fd_sc_hd__xnor2_1 _16219_ (.A(_09192_),
    .B(_09311_),
    .Y(_09312_));
 sky130_fd_sc_hd__xor2_2 _16220_ (.A(_09307_),
    .B(_09312_),
    .X(_09313_));
 sky130_fd_sc_hd__nand2_1 _16221_ (.A(_08466_),
    .B(_09184_),
    .Y(_09314_));
 sky130_fd_sc_hd__clkbuf_4 _16222_ (.A(_09053_),
    .X(_09315_));
 sky130_fd_sc_hd__o22ai_1 _16223_ (.A1(_08581_),
    .A2(_09315_),
    .B1(_09195_),
    .B2(_08461_),
    .Y(_09316_));
 sky130_fd_sc_hd__a31o_1 _16224_ (.A1(_08733_),
    .A2(_09314_),
    .A3(_09316_),
    .B1(_09193_),
    .X(_09317_));
 sky130_fd_sc_hd__xor2_2 _16225_ (.A(_09313_),
    .B(_09317_),
    .X(_09318_));
 sky130_fd_sc_hd__xnor2_2 _16226_ (.A(_09305_),
    .B(_09318_),
    .Y(_09319_));
 sky130_fd_sc_hd__and3_1 _16227_ (.A(_09197_),
    .B(_09198_),
    .C(_09201_),
    .X(_09320_));
 sky130_fd_sc_hd__a21oi_1 _16228_ (.A1(_09183_),
    .A2(_09202_),
    .B1(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__xor2_1 _16229_ (.A(_09319_),
    .B(_09321_),
    .X(_09322_));
 sky130_fd_sc_hd__xnor2_1 _16230_ (.A(_09301_),
    .B(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__and2b_1 _16231_ (.A_N(_09203_),
    .B(_09205_),
    .X(_09324_));
 sky130_fd_sc_hd__a21oi_1 _16232_ (.A1(_09175_),
    .A2(_09206_),
    .B1(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__nor2_1 _16233_ (.A(_09323_),
    .B(_09325_),
    .Y(_09326_));
 sky130_fd_sc_hd__and2_1 _16234_ (.A(_09323_),
    .B(_09325_),
    .X(_09327_));
 sky130_fd_sc_hd__nor2_1 _16235_ (.A(_09326_),
    .B(_09327_),
    .Y(_09328_));
 sky130_fd_sc_hd__xnor2_2 _16236_ (.A(_09288_),
    .B(_09328_),
    .Y(_09329_));
 sky130_fd_sc_hd__nor2_1 _16237_ (.A(_09207_),
    .B(_09209_),
    .Y(_09330_));
 sky130_fd_sc_hd__a21oi_1 _16238_ (.A1(_09165_),
    .A2(_09210_),
    .B1(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__xor2_1 _16239_ (.A(_09329_),
    .B(_09331_),
    .X(_09332_));
 sky130_fd_sc_hd__xnor2_1 _16240_ (.A(_09267_),
    .B(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__a21oi_1 _16241_ (.A1(_09143_),
    .A2(_09216_),
    .B1(_09214_),
    .Y(_09334_));
 sky130_fd_sc_hd__nor2_1 _16242_ (.A(_09333_),
    .B(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__and2_1 _16243_ (.A(_09333_),
    .B(_09334_),
    .X(_09336_));
 sky130_fd_sc_hd__nor2_1 _16244_ (.A(_09335_),
    .B(_09336_),
    .Y(_09337_));
 sky130_fd_sc_hd__xnor2_1 _16245_ (.A(_09239_),
    .B(_09337_),
    .Y(_09338_));
 sky130_fd_sc_hd__a21oi_1 _16246_ (.A1(_09086_),
    .A2(_09220_),
    .B1(_09219_),
    .Y(_09339_));
 sky130_fd_sc_hd__or2_2 _16247_ (.A(_09338_),
    .B(_09339_),
    .X(_09340_));
 sky130_fd_sc_hd__nand2_1 _16248_ (.A(_09338_),
    .B(_09339_),
    .Y(_09341_));
 sky130_fd_sc_hd__or4bb_1 _16249_ (.A(_09222_),
    .B(_09224_),
    .C_N(_09340_),
    .D_N(_09341_),
    .X(_09342_));
 sky130_fd_sc_hd__a2bb2o_1 _16250_ (.A1_N(_09222_),
    .A2_N(_09224_),
    .B1(_09340_),
    .B2(_09341_),
    .X(_09343_));
 sky130_fd_sc_hd__and2_2 _16251_ (.A(_09342_),
    .B(_09343_),
    .X(_09344_));
 sky130_fd_sc_hd__a21oi_1 _16252_ (.A1(_09126_),
    .A2(_09098_),
    .B1(_09225_),
    .Y(_09345_));
 sky130_fd_sc_hd__a31o_4 _16253_ (.A1(_09000_),
    .A2(_09100_),
    .A3(_09226_),
    .B1(_09345_),
    .X(_09346_));
 sky130_fd_sc_hd__xor2_4 _16254_ (.A(_09344_),
    .B(_09346_),
    .X(_09347_));
 sky130_fd_sc_hd__mux2_1 _16255_ (.A0(\rbzero.debug_overlay.playerY[-4] ),
    .A1(\rbzero.debug_overlay.playerX[-4] ),
    .S(_08138_),
    .X(_09348_));
 sky130_fd_sc_hd__xnor2_1 _16256_ (.A(_09347_),
    .B(_09348_),
    .Y(_09349_));
 sky130_fd_sc_hd__a21oi_1 _16257_ (.A1(_09238_),
    .A2(_09232_),
    .B1(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__and3_1 _16258_ (.A(_09238_),
    .B(_09232_),
    .C(_09349_),
    .X(_09351_));
 sky130_fd_sc_hd__nor2_1 _16259_ (.A(_09350_),
    .B(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__xnor2_1 _16260_ (.A(_09121_),
    .B(_09352_),
    .Y(_09353_));
 sky130_fd_sc_hd__nand2_1 _16261_ (.A(_08145_),
    .B(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__o211a_1 _16262_ (.A1(\rbzero.texu_hot[2] ),
    .A2(_08145_),
    .B1(_09354_),
    .C1(_08085_),
    .X(_00468_));
 sky130_fd_sc_hd__a21boi_4 _16263_ (.A1(_09344_),
    .A2(_09346_),
    .B1_N(_09342_),
    .Y(_09355_));
 sky130_fd_sc_hd__a21o_1 _16264_ (.A1(_09162_),
    .A2(_09240_),
    .B1(_09264_),
    .X(_09356_));
 sky130_fd_sc_hd__o21ai_1 _16265_ (.A1(_09265_),
    .A2(_09266_),
    .B1(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__nand2_1 _16266_ (.A(_09244_),
    .B(_09263_),
    .Y(_09358_));
 sky130_fd_sc_hd__o21ai_1 _16267_ (.A1(_09260_),
    .A2(_09262_),
    .B1(_09358_),
    .Y(_09359_));
 sky130_fd_sc_hd__or2b_1 _16268_ (.A(_09287_),
    .B_N(_09268_),
    .X(_09360_));
 sky130_fd_sc_hd__a21bo_1 _16269_ (.A1(_09270_),
    .A2(_09286_),
    .B1_N(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__nand2_4 _16270_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_08475_),
    .Y(_09362_));
 sky130_fd_sc_hd__buf_4 _16271_ (.A(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__nor2_1 _16272_ (.A(_08304_),
    .B(_09363_),
    .Y(_09364_));
 sky130_fd_sc_hd__nor2_1 _16273_ (.A(_08304_),
    .B(_09243_),
    .Y(_09365_));
 sky130_fd_sc_hd__o21ba_1 _16274_ (.A1(_08616_),
    .A2(_09363_),
    .B1_N(_09365_),
    .X(_09366_));
 sky130_fd_sc_hd__a21oi_1 _16275_ (.A1(_09244_),
    .A2(_09364_),
    .B1(_09366_),
    .Y(_09367_));
 sky130_fd_sc_hd__a21bo_1 _16276_ (.A1(_09248_),
    .A2(_09249_),
    .B1_N(_09251_),
    .X(_09368_));
 sky130_fd_sc_hd__or3_1 _16277_ (.A(_09005_),
    .B(_08553_),
    .C(_09273_),
    .X(_09369_));
 sky130_fd_sc_hd__nor2_1 _16278_ (.A(_08296_),
    .B(_09076_),
    .Y(_09370_));
 sky130_fd_sc_hd__nor2_1 _16279_ (.A(_08274_),
    .B(_08617_),
    .Y(_09371_));
 sky130_fd_sc_hd__xnor2_1 _16280_ (.A(_09370_),
    .B(_09371_),
    .Y(_09372_));
 sky130_fd_sc_hd__or3_1 _16281_ (.A(_08335_),
    .B(_09131_),
    .C(_09372_),
    .X(_09373_));
 sky130_fd_sc_hd__o21ai_1 _16282_ (.A1(_09008_),
    .A2(_09131_),
    .B1(_09372_),
    .Y(_09374_));
 sky130_fd_sc_hd__nand2_1 _16283_ (.A(_09373_),
    .B(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__a21o_1 _16284_ (.A1(_09271_),
    .A2(_09369_),
    .B1(_09375_),
    .X(_09376_));
 sky130_fd_sc_hd__nand3_1 _16285_ (.A(_09271_),
    .B(_09369_),
    .C(_09375_),
    .Y(_09377_));
 sky130_fd_sc_hd__nand2_1 _16286_ (.A(_09376_),
    .B(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__xor2_1 _16287_ (.A(_09368_),
    .B(_09378_),
    .X(_09379_));
 sky130_fd_sc_hd__o21a_1 _16288_ (.A1(_09247_),
    .A2(_09259_),
    .B1(_09257_),
    .X(_09380_));
 sky130_fd_sc_hd__xor2_1 _16289_ (.A(_09379_),
    .B(_09380_),
    .X(_09381_));
 sky130_fd_sc_hd__xor2_1 _16290_ (.A(_09367_),
    .B(_09381_),
    .X(_09382_));
 sky130_fd_sc_hd__xnor2_1 _16291_ (.A(_09361_),
    .B(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__xnor2_1 _16292_ (.A(_09359_),
    .B(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__o21ai_1 _16293_ (.A1(_09280_),
    .A2(_09282_),
    .B1(_09284_),
    .Y(_09385_));
 sky130_fd_sc_hd__a21bo_1 _16294_ (.A1(_09289_),
    .A2(_09299_),
    .B1_N(_09298_),
    .X(_09386_));
 sky130_fd_sc_hd__o22ai_1 _16295_ (.A1(_08151_),
    .A2(_08734_),
    .B1(_08731_),
    .B2(_08166_),
    .Y(_09387_));
 sky130_fd_sc_hd__or4_1 _16296_ (.A(_08151_),
    .B(_08165_),
    .C(_08734_),
    .D(_08731_),
    .X(_09388_));
 sky130_fd_sc_hd__nand2_1 _16297_ (.A(_09387_),
    .B(_09388_),
    .Y(_09389_));
 sky130_fd_sc_hd__or3_1 _16298_ (.A(_09146_),
    .B(_08553_),
    .C(_09389_),
    .X(_09390_));
 sky130_fd_sc_hd__o21ai_1 _16299_ (.A1(_09146_),
    .A2(_08620_),
    .B1(_09389_),
    .Y(_09391_));
 sky130_fd_sc_hd__and2_1 _16300_ (.A(_09390_),
    .B(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__nor2_2 _16301_ (.A(_08813_),
    .B(_08409_),
    .Y(_09393_));
 sky130_fd_sc_hd__xnor2_1 _16302_ (.A(_09276_),
    .B(_09393_),
    .Y(_09394_));
 sky130_fd_sc_hd__or2_1 _16303_ (.A(_08368_),
    .B(_08535_),
    .X(_09395_));
 sky130_fd_sc_hd__xnor2_1 _16304_ (.A(_09394_),
    .B(_09395_),
    .Y(_09396_));
 sky130_fd_sc_hd__clkbuf_4 _16305_ (.A(_08535_),
    .X(_09397_));
 sky130_fd_sc_hd__nand2_1 _16306_ (.A(_09152_),
    .B(_09276_),
    .Y(_09398_));
 sky130_fd_sc_hd__o31a_1 _16307_ (.A1(_08370_),
    .A2(_09397_),
    .A3(_09277_),
    .B1(_09398_),
    .X(_09399_));
 sky130_fd_sc_hd__nor2_1 _16308_ (.A(_09396_),
    .B(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__and2_1 _16309_ (.A(_09396_),
    .B(_09399_),
    .X(_09401_));
 sky130_fd_sc_hd__nor2_1 _16310_ (.A(_09400_),
    .B(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__xor2_1 _16311_ (.A(_09392_),
    .B(_09402_),
    .X(_09403_));
 sky130_fd_sc_hd__xnor2_1 _16312_ (.A(_09386_),
    .B(_09403_),
    .Y(_09404_));
 sky130_fd_sc_hd__xnor2_1 _16313_ (.A(_09385_),
    .B(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__clkbuf_4 _16314_ (.A(_08373_),
    .X(_09406_));
 sky130_fd_sc_hd__nand2_1 _16315_ (.A(_09170_),
    .B(_09293_),
    .Y(_09407_));
 sky130_fd_sc_hd__o31ai_1 _16316_ (.A1(_09406_),
    .A2(_08409_),
    .A3(_09294_),
    .B1(_09407_),
    .Y(_09408_));
 sky130_fd_sc_hd__a22o_1 _16317_ (.A1(_09290_),
    .A2(_09303_),
    .B1(_09304_),
    .B2(_09302_),
    .X(_09409_));
 sky130_fd_sc_hd__nor2_1 _16318_ (.A(_08369_),
    .B(_09037_),
    .Y(_09410_));
 sky130_fd_sc_hd__xnor2_1 _16319_ (.A(_09293_),
    .B(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__nor2_1 _16320_ (.A(_08373_),
    .B(_08497_),
    .Y(_09412_));
 sky130_fd_sc_hd__xnor2_1 _16321_ (.A(_09411_),
    .B(_09412_),
    .Y(_09413_));
 sky130_fd_sc_hd__xnor2_1 _16322_ (.A(_09409_),
    .B(_09413_),
    .Y(_09414_));
 sky130_fd_sc_hd__xnor2_1 _16323_ (.A(_09408_),
    .B(_09414_),
    .Y(_09415_));
 sky130_fd_sc_hd__a21oi_1 _16324_ (.A1(_09044_),
    .A2(_09046_),
    .B1(_08434_),
    .Y(_09416_));
 sky130_fd_sc_hd__a21o_1 _16325_ (.A1(_08466_),
    .A2(_09184_),
    .B1(_08910_),
    .X(_09417_));
 sky130_fd_sc_hd__a21oi_1 _16326_ (.A1(_09315_),
    .A2(_09306_),
    .B1(_08431_),
    .Y(_09418_));
 sky130_fd_sc_hd__xnor2_1 _16327_ (.A(_09417_),
    .B(_09418_),
    .Y(_09419_));
 sky130_fd_sc_hd__xor2_1 _16328_ (.A(_09416_),
    .B(_09419_),
    .X(_09420_));
 sky130_fd_sc_hd__nand2_2 _16329_ (.A(\rbzero.wall_tracer.stepDistX[6] ),
    .B(_09045_),
    .Y(_09421_));
 sky130_fd_sc_hd__and2_1 _16330_ (.A(_09195_),
    .B(_09421_),
    .X(_09422_));
 sky130_fd_sc_hd__inv_2 _16331_ (.A(_08026_),
    .Y(_09423_));
 sky130_fd_sc_hd__o41a_1 _16332_ (.A1(_08012_),
    .A2(_08023_),
    .A3(_08450_),
    .A4(_09188_),
    .B1(_08027_),
    .X(_09424_));
 sky130_fd_sc_hd__a211o_1 _16333_ (.A1(_09423_),
    .A2(_09308_),
    .B1(_09424_),
    .C1(_08144_),
    .X(_09425_));
 sky130_fd_sc_hd__a22o_2 _16334_ (.A1(\rbzero.wall_tracer.stepDistY[8] ),
    .A2(_08405_),
    .B1(_09190_),
    .B2(_09425_),
    .X(_09426_));
 sky130_fd_sc_hd__nand3_1 _16335_ (.A(_08471_),
    .B(_09311_),
    .C(_09426_),
    .Y(_09427_));
 sky130_fd_sc_hd__and3_1 _16336_ (.A(\rbzero.wall_tracer.visualWallDist[-10] ),
    .B(_08149_),
    .C(_09310_),
    .X(_09428_));
 sky130_fd_sc_hd__a21o_1 _16337_ (.A1(_08484_),
    .A2(_09426_),
    .B1(_09428_),
    .X(_09429_));
 sky130_fd_sc_hd__or4bb_1 _16338_ (.A(_08441_),
    .B(_09422_),
    .C_N(_09427_),
    .D_N(_09429_),
    .X(_09430_));
 sky130_fd_sc_hd__a2bb2o_1 _16339_ (.A1_N(_08441_),
    .A2_N(_09422_),
    .B1(_09427_),
    .B2(_09429_),
    .X(_09431_));
 sky130_fd_sc_hd__and3_1 _16340_ (.A(\rbzero.trace_state[0] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .C(_08338_),
    .X(_09432_));
 sky130_fd_sc_hd__o21ai_4 _16341_ (.A1(_09432_),
    .A2(_09310_),
    .B1(_06263_),
    .Y(_09433_));
 sky130_fd_sc_hd__or3_1 _16342_ (.A(_08461_),
    .B(_09192_),
    .C(_09433_),
    .X(_09434_));
 sky130_fd_sc_hd__a21bo_1 _16343_ (.A1(_09307_),
    .A2(_09312_),
    .B1_N(_09434_),
    .X(_09435_));
 sky130_fd_sc_hd__nand3_1 _16344_ (.A(_09430_),
    .B(_09431_),
    .C(_09435_),
    .Y(_09436_));
 sky130_fd_sc_hd__a21o_1 _16345_ (.A1(_09430_),
    .A2(_09431_),
    .B1(_09435_),
    .X(_09437_));
 sky130_fd_sc_hd__nand3_1 _16346_ (.A(_09420_),
    .B(_09436_),
    .C(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__a21o_1 _16347_ (.A1(_09436_),
    .A2(_09437_),
    .B1(_09420_),
    .X(_09439_));
 sky130_fd_sc_hd__and2_1 _16348_ (.A(_09313_),
    .B(_09317_),
    .X(_09440_));
 sky130_fd_sc_hd__a21o_1 _16349_ (.A1(_09305_),
    .A2(_09318_),
    .B1(_09440_),
    .X(_09441_));
 sky130_fd_sc_hd__nand3_1 _16350_ (.A(_09438_),
    .B(_09439_),
    .C(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__a21o_1 _16351_ (.A1(_09438_),
    .A2(_09439_),
    .B1(_09441_),
    .X(_09443_));
 sky130_fd_sc_hd__and3_1 _16352_ (.A(_09415_),
    .B(_09442_),
    .C(_09443_),
    .X(_09444_));
 sky130_fd_sc_hd__a21oi_1 _16353_ (.A1(_09442_),
    .A2(_09443_),
    .B1(_09415_),
    .Y(_09445_));
 sky130_fd_sc_hd__or2_1 _16354_ (.A(_09444_),
    .B(_09445_),
    .X(_09446_));
 sky130_fd_sc_hd__nor2_1 _16355_ (.A(_09319_),
    .B(_09321_),
    .Y(_09447_));
 sky130_fd_sc_hd__a21oi_1 _16356_ (.A1(_09301_),
    .A2(_09322_),
    .B1(_09447_),
    .Y(_09448_));
 sky130_fd_sc_hd__nor2_1 _16357_ (.A(_09446_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__nand2_1 _16358_ (.A(_09446_),
    .B(_09448_),
    .Y(_09450_));
 sky130_fd_sc_hd__and2b_1 _16359_ (.A_N(_09449_),
    .B(_09450_),
    .X(_09451_));
 sky130_fd_sc_hd__xnor2_1 _16360_ (.A(_09405_),
    .B(_09451_),
    .Y(_09452_));
 sky130_fd_sc_hd__a21oi_1 _16361_ (.A1(_09288_),
    .A2(_09328_),
    .B1(_09326_),
    .Y(_09453_));
 sky130_fd_sc_hd__nor2_1 _16362_ (.A(_09452_),
    .B(_09453_),
    .Y(_09454_));
 sky130_fd_sc_hd__and2_1 _16363_ (.A(_09452_),
    .B(_09453_),
    .X(_09455_));
 sky130_fd_sc_hd__nor2_1 _16364_ (.A(_09454_),
    .B(_09455_),
    .Y(_09456_));
 sky130_fd_sc_hd__xnor2_1 _16365_ (.A(_09384_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__nor2_1 _16366_ (.A(_09329_),
    .B(_09331_),
    .Y(_09458_));
 sky130_fd_sc_hd__a21oi_1 _16367_ (.A1(_09267_),
    .A2(_09332_),
    .B1(_09458_),
    .Y(_09459_));
 sky130_fd_sc_hd__xnor2_1 _16368_ (.A(_09457_),
    .B(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__xor2_1 _16369_ (.A(_09357_),
    .B(_09460_),
    .X(_09461_));
 sky130_fd_sc_hd__a21oi_1 _16370_ (.A1(_09239_),
    .A2(_09337_),
    .B1(_09335_),
    .Y(_09462_));
 sky130_fd_sc_hd__nor2_1 _16371_ (.A(_09461_),
    .B(_09462_),
    .Y(_09463_));
 sky130_fd_sc_hd__and2_1 _16372_ (.A(_09461_),
    .B(_09462_),
    .X(_09464_));
 sky130_fd_sc_hd__or2_2 _16373_ (.A(_09463_),
    .B(_09464_),
    .X(_09465_));
 sky130_fd_sc_hd__xor2_4 _16374_ (.A(_09340_),
    .B(_09465_),
    .X(_09466_));
 sky130_fd_sc_hd__xor2_4 _16375_ (.A(_09355_),
    .B(_09466_),
    .X(_09467_));
 sky130_fd_sc_hd__clkinv_2 _16376_ (.A(\rbzero.debug_overlay.playerX[-3] ),
    .Y(_09468_));
 sky130_fd_sc_hd__mux2_1 _16377_ (.A0(_04686_),
    .A1(_09468_),
    .S(_08138_),
    .X(_09469_));
 sky130_fd_sc_hd__nor2_1 _16378_ (.A(_09467_),
    .B(_09469_),
    .Y(_09470_));
 sky130_fd_sc_hd__and2_1 _16379_ (.A(_09467_),
    .B(_09469_),
    .X(_09471_));
 sky130_fd_sc_hd__or2_1 _16380_ (.A(_09470_),
    .B(_09471_),
    .X(_09472_));
 sky130_fd_sc_hd__a21oi_1 _16381_ (.A1(_09347_),
    .A2(_09348_),
    .B1(_09350_),
    .Y(_09473_));
 sky130_fd_sc_hd__xnor2_1 _16382_ (.A(_09472_),
    .B(_09473_),
    .Y(_09474_));
 sky130_fd_sc_hd__o21ai_1 _16383_ (.A1(_09121_),
    .A2(_09474_),
    .B1(_08145_),
    .Y(_09475_));
 sky130_fd_sc_hd__a21o_1 _16384_ (.A1(_09121_),
    .A2(_09474_),
    .B1(_09475_),
    .X(_09476_));
 sky130_fd_sc_hd__o211a_1 _16385_ (.A1(\rbzero.texu_hot[3] ),
    .A2(_08145_),
    .B1(_09476_),
    .C1(_08085_),
    .X(_00469_));
 sky130_fd_sc_hd__o21ba_1 _16386_ (.A1(_09472_),
    .A2(_09473_),
    .B1_N(_09470_),
    .X(_09477_));
 sky130_fd_sc_hd__a21oi_1 _16387_ (.A1(_09340_),
    .A2(_09342_),
    .B1(_09465_),
    .Y(_09478_));
 sky130_fd_sc_hd__a31oi_4 _16388_ (.A1(_09344_),
    .A2(_09346_),
    .A3(_09466_),
    .B1(_09478_),
    .Y(_09479_));
 sky130_fd_sc_hd__or2_1 _16389_ (.A(_09457_),
    .B(_09459_),
    .X(_09480_));
 sky130_fd_sc_hd__or2b_1 _16390_ (.A(_09460_),
    .B_N(_09357_),
    .X(_09481_));
 sky130_fd_sc_hd__or2b_1 _16391_ (.A(_09383_),
    .B_N(_09359_),
    .X(_09482_));
 sky130_fd_sc_hd__a21bo_1 _16392_ (.A1(_09361_),
    .A2(_09382_),
    .B1_N(_09482_),
    .X(_09483_));
 sky130_fd_sc_hd__a2bb2o_1 _16393_ (.A1_N(_09379_),
    .A2_N(_09380_),
    .B1(_09381_),
    .B2(_09367_),
    .X(_09484_));
 sky130_fd_sc_hd__nand2_1 _16394_ (.A(_09386_),
    .B(_09403_),
    .Y(_09485_));
 sky130_fd_sc_hd__or2b_1 _16395_ (.A(_09404_),
    .B_N(_09385_),
    .X(_09486_));
 sky130_fd_sc_hd__nand2_1 _16396_ (.A(_09244_),
    .B(_09364_),
    .Y(_09487_));
 sky130_fd_sc_hd__nor2_1 _16397_ (.A(_09008_),
    .B(_09242_),
    .Y(_09488_));
 sky130_fd_sc_hd__xnor2_1 _16398_ (.A(_09364_),
    .B(_09488_),
    .Y(_09489_));
 sky130_fd_sc_hd__nand2_2 _16399_ (.A(\rbzero.wall_tracer.visualWallDist[9] ),
    .B(_08475_),
    .Y(_09490_));
 sky130_fd_sc_hd__clkbuf_4 _16400_ (.A(_09490_),
    .X(_09491_));
 sky130_fd_sc_hd__nor3_1 _16401_ (.A(_08616_),
    .B(_09489_),
    .C(_09491_),
    .Y(_09492_));
 sky130_fd_sc_hd__o21a_1 _16402_ (.A1(_08616_),
    .A2(_09491_),
    .B1(_09489_),
    .X(_09493_));
 sky130_fd_sc_hd__nor2_1 _16403_ (.A(_09492_),
    .B(_09493_),
    .Y(_09494_));
 sky130_fd_sc_hd__xnor2_1 _16404_ (.A(_09487_),
    .B(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__or2b_1 _16405_ (.A(_09378_),
    .B_N(_09368_),
    .X(_09496_));
 sky130_fd_sc_hd__a21bo_1 _16406_ (.A1(_09370_),
    .A2(_09371_),
    .B1_N(_09373_),
    .X(_09497_));
 sky130_fd_sc_hd__nor2_2 _16407_ (.A(_08952_),
    .B(_09131_),
    .Y(_09498_));
 sky130_fd_sc_hd__nor2_1 _16408_ (.A(_08847_),
    .B(_09076_),
    .Y(_09499_));
 sky130_fd_sc_hd__o22a_1 _16409_ (.A1(_08847_),
    .A2(_08617_),
    .B1(_09076_),
    .B2(_08274_),
    .X(_09500_));
 sky130_fd_sc_hd__a21oi_1 _16410_ (.A1(_09371_),
    .A2(_09499_),
    .B1(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__xnor2_1 _16411_ (.A(_09498_),
    .B(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__a21oi_1 _16412_ (.A1(_09388_),
    .A2(_09390_),
    .B1(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__and3_1 _16413_ (.A(_09388_),
    .B(_09390_),
    .C(_09502_),
    .X(_09504_));
 sky130_fd_sc_hd__nor2_1 _16414_ (.A(_09503_),
    .B(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__xnor2_1 _16415_ (.A(_09497_),
    .B(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__a21oi_1 _16416_ (.A1(_09376_),
    .A2(_09496_),
    .B1(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__and3_1 _16417_ (.A(_09376_),
    .B(_09496_),
    .C(_09506_),
    .X(_09508_));
 sky130_fd_sc_hd__nor2_1 _16418_ (.A(_09507_),
    .B(_09508_),
    .Y(_09509_));
 sky130_fd_sc_hd__xnor2_1 _16419_ (.A(_09495_),
    .B(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__a21o_1 _16420_ (.A1(_09485_),
    .A2(_09486_),
    .B1(_09510_),
    .X(_09511_));
 sky130_fd_sc_hd__nand3_1 _16421_ (.A(_09485_),
    .B(_09486_),
    .C(_09510_),
    .Y(_09512_));
 sky130_fd_sc_hd__nand2_1 _16422_ (.A(_09511_),
    .B(_09512_),
    .Y(_09513_));
 sky130_fd_sc_hd__xnor2_1 _16423_ (.A(_09484_),
    .B(_09513_),
    .Y(_09514_));
 sky130_fd_sc_hd__a21o_1 _16424_ (.A1(_09392_),
    .A2(_09402_),
    .B1(_09400_),
    .X(_09515_));
 sky130_fd_sc_hd__or2_1 _16425_ (.A(_09409_),
    .B(_09413_),
    .X(_09516_));
 sky130_fd_sc_hd__and2_1 _16426_ (.A(_09409_),
    .B(_09413_),
    .X(_09517_));
 sky130_fd_sc_hd__a21o_1 _16427_ (.A1(_09408_),
    .A2(_09516_),
    .B1(_09517_),
    .X(_09518_));
 sky130_fd_sc_hd__clkbuf_4 _16428_ (.A(_08666_),
    .X(_09519_));
 sky130_fd_sc_hd__clkbuf_4 _16429_ (.A(_08734_),
    .X(_09520_));
 sky130_fd_sc_hd__o22ai_1 _16430_ (.A1(_08152_),
    .A2(_09519_),
    .B1(_09520_),
    .B2(_08166_),
    .Y(_09521_));
 sky130_fd_sc_hd__or2_1 _16431_ (.A(_08166_),
    .B(_08666_),
    .X(_09522_));
 sky130_fd_sc_hd__or3_1 _16432_ (.A(_08152_),
    .B(_09520_),
    .C(_09522_),
    .X(_09523_));
 sky130_fd_sc_hd__nand2_1 _16433_ (.A(_09521_),
    .B(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__buf_2 _16434_ (.A(_08731_),
    .X(_09525_));
 sky130_fd_sc_hd__nor2_1 _16435_ (.A(_09525_),
    .B(_08620_),
    .Y(_09526_));
 sky130_fd_sc_hd__xnor2_1 _16436_ (.A(_09524_),
    .B(_09526_),
    .Y(_09527_));
 sky130_fd_sc_hd__clkbuf_4 _16437_ (.A(_08327_),
    .X(_09528_));
 sky130_fd_sc_hd__nor2_2 _16438_ (.A(_09528_),
    .B(_08497_),
    .Y(_09529_));
 sky130_fd_sc_hd__o22a_1 _16439_ (.A1(_08813_),
    .A2(_08497_),
    .B1(_08409_),
    .B2(_09528_),
    .X(_09530_));
 sky130_fd_sc_hd__a21oi_1 _16440_ (.A1(_09393_),
    .A2(_09529_),
    .B1(_09530_),
    .Y(_09531_));
 sky130_fd_sc_hd__nor2_1 _16441_ (.A(_09397_),
    .B(_08384_),
    .Y(_09532_));
 sky130_fd_sc_hd__xnor2_1 _16442_ (.A(_09531_),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__nand2_1 _16443_ (.A(_09276_),
    .B(_09393_),
    .Y(_09534_));
 sky130_fd_sc_hd__o31a_1 _16444_ (.A1(_08368_),
    .A2(_09397_),
    .A3(_09394_),
    .B1(_09534_),
    .X(_09535_));
 sky130_fd_sc_hd__nor2_1 _16445_ (.A(_09533_),
    .B(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__nand2_1 _16446_ (.A(_09533_),
    .B(_09535_),
    .Y(_09537_));
 sky130_fd_sc_hd__and2b_1 _16447_ (.A_N(_09536_),
    .B(_09537_),
    .X(_09538_));
 sky130_fd_sc_hd__xnor2_1 _16448_ (.A(_09527_),
    .B(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__xor2_1 _16449_ (.A(_09518_),
    .B(_09539_),
    .X(_09540_));
 sky130_fd_sc_hd__xnor2_1 _16450_ (.A(_09515_),
    .B(_09540_),
    .Y(_09541_));
 sky130_fd_sc_hd__clkbuf_4 _16451_ (.A(_09406_),
    .X(_09542_));
 sky130_fd_sc_hd__or3_1 _16452_ (.A(_09542_),
    .B(_08497_),
    .C(_09411_),
    .X(_09543_));
 sky130_fd_sc_hd__a21bo_1 _16453_ (.A1(_09293_),
    .A2(_09410_),
    .B1_N(_09543_),
    .X(_09544_));
 sky130_fd_sc_hd__a21oi_2 _16454_ (.A1(_09053_),
    .A2(_09306_),
    .B1(_08910_),
    .Y(_09545_));
 sky130_fd_sc_hd__a22o_1 _16455_ (.A1(_09303_),
    .A2(_09545_),
    .B1(_09419_),
    .B2(_09416_),
    .X(_09546_));
 sky130_fd_sc_hd__nor2_1 _16456_ (.A(_08516_),
    .B(_09037_),
    .Y(_09547_));
 sky130_fd_sc_hd__a21oi_1 _16457_ (.A1(_09044_),
    .A2(_09046_),
    .B1(_08369_),
    .Y(_09548_));
 sky130_fd_sc_hd__xnor2_1 _16458_ (.A(_09547_),
    .B(_09548_),
    .Y(_09549_));
 sky130_fd_sc_hd__or3_1 _16459_ (.A(_09406_),
    .B(_09176_),
    .C(_09549_),
    .X(_09550_));
 sky130_fd_sc_hd__o21ai_1 _16460_ (.A1(_09406_),
    .A2(_09176_),
    .B1(_09549_),
    .Y(_09551_));
 sky130_fd_sc_hd__and2_1 _16461_ (.A(_09550_),
    .B(_09551_),
    .X(_09552_));
 sky130_fd_sc_hd__xor2_2 _16462_ (.A(_09546_),
    .B(_09552_),
    .X(_09553_));
 sky130_fd_sc_hd__xor2_2 _16463_ (.A(_09544_),
    .B(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__a21oi_1 _16464_ (.A1(_09195_),
    .A2(_09421_),
    .B1(_08431_),
    .Y(_09555_));
 sky130_fd_sc_hd__xnor2_1 _16465_ (.A(_09545_),
    .B(_09555_),
    .Y(_09556_));
 sky130_fd_sc_hd__nor2_1 _16466_ (.A(_08434_),
    .B(_09186_),
    .Y(_09557_));
 sky130_fd_sc_hd__xnor2_2 _16467_ (.A(_09556_),
    .B(_09557_),
    .Y(_09558_));
 sky130_fd_sc_hd__a21boi_4 _16468_ (.A1(\rbzero.wall_tracer.stepDistX[7] ),
    .A2(_09045_),
    .B1_N(_09433_),
    .Y(_09559_));
 sky130_fd_sc_hd__clkbuf_4 _16469_ (.A(_09559_),
    .X(_09560_));
 sky130_fd_sc_hd__nor2_1 _16470_ (.A(_08950_),
    .B(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__nand2_1 _16471_ (.A(_08471_),
    .B(_09426_),
    .Y(_09562_));
 sky130_fd_sc_hd__or4_1 _16472_ (.A(_08011_),
    .B(_08023_),
    .C(_08449_),
    .D(_09188_),
    .X(_09563_));
 sky130_fd_sc_hd__or3_1 _16473_ (.A(_08027_),
    .B(_08029_),
    .C(_09563_),
    .X(_09564_));
 sky130_fd_sc_hd__o21ai_1 _16474_ (.A1(_08027_),
    .A2(_09563_),
    .B1(_08029_),
    .Y(_09565_));
 sky130_fd_sc_hd__a31o_1 _16475_ (.A1(_08148_),
    .A2(_09564_),
    .A3(_09565_),
    .B1(_08454_),
    .X(_09566_));
 sky130_fd_sc_hd__or3_2 _16476_ (.A(_08039_),
    .B(_08338_),
    .C(_09566_),
    .X(_09567_));
 sky130_fd_sc_hd__xor2_2 _16477_ (.A(_09562_),
    .B(_09567_),
    .X(_09568_));
 sky130_fd_sc_hd__xnor2_2 _16478_ (.A(_09561_),
    .B(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__nand2_1 _16479_ (.A(_09427_),
    .B(_09430_),
    .Y(_09570_));
 sky130_fd_sc_hd__xnor2_2 _16480_ (.A(_09569_),
    .B(_09570_),
    .Y(_09571_));
 sky130_fd_sc_hd__xnor2_2 _16481_ (.A(_09558_),
    .B(_09571_),
    .Y(_09572_));
 sky130_fd_sc_hd__and2_1 _16482_ (.A(_09436_),
    .B(_09438_),
    .X(_09573_));
 sky130_fd_sc_hd__xor2_2 _16483_ (.A(_09572_),
    .B(_09573_),
    .X(_09574_));
 sky130_fd_sc_hd__xnor2_2 _16484_ (.A(_09554_),
    .B(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__a21boi_2 _16485_ (.A1(_09415_),
    .A2(_09443_),
    .B1_N(_09442_),
    .Y(_09576_));
 sky130_fd_sc_hd__xor2_1 _16486_ (.A(_09575_),
    .B(_09576_),
    .X(_09577_));
 sky130_fd_sc_hd__xnor2_1 _16487_ (.A(_09541_),
    .B(_09577_),
    .Y(_09578_));
 sky130_fd_sc_hd__a21oi_1 _16488_ (.A1(_09405_),
    .A2(_09451_),
    .B1(_09449_),
    .Y(_09579_));
 sky130_fd_sc_hd__nor2_1 _16489_ (.A(_09578_),
    .B(_09579_),
    .Y(_09580_));
 sky130_fd_sc_hd__nand2_1 _16490_ (.A(_09578_),
    .B(_09579_),
    .Y(_09581_));
 sky130_fd_sc_hd__and2b_1 _16491_ (.A_N(_09580_),
    .B(_09581_),
    .X(_09582_));
 sky130_fd_sc_hd__xnor2_1 _16492_ (.A(_09514_),
    .B(_09582_),
    .Y(_09583_));
 sky130_fd_sc_hd__a21oi_1 _16493_ (.A1(_09384_),
    .A2(_09456_),
    .B1(_09454_),
    .Y(_09584_));
 sky130_fd_sc_hd__xor2_1 _16494_ (.A(_09583_),
    .B(_09584_),
    .X(_09585_));
 sky130_fd_sc_hd__xnor2_1 _16495_ (.A(_09483_),
    .B(_09585_),
    .Y(_09586_));
 sky130_fd_sc_hd__a21o_2 _16496_ (.A1(_09480_),
    .A2(_09481_),
    .B1(_09586_),
    .X(_09587_));
 sky130_fd_sc_hd__nand3_1 _16497_ (.A(_09480_),
    .B(_09481_),
    .C(_09586_),
    .Y(_09588_));
 sky130_fd_sc_hd__and2_1 _16498_ (.A(_09587_),
    .B(_09588_),
    .X(_09589_));
 sky130_fd_sc_hd__nand2_1 _16499_ (.A(_09463_),
    .B(_09589_),
    .Y(_09590_));
 sky130_fd_sc_hd__or2_1 _16500_ (.A(_09463_),
    .B(_09589_),
    .X(_09591_));
 sky130_fd_sc_hd__nand2_2 _16501_ (.A(_09590_),
    .B(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__xor2_4 _16502_ (.A(_09479_),
    .B(_09592_),
    .X(_09593_));
 sky130_fd_sc_hd__mux2_1 _16503_ (.A0(\rbzero.debug_overlay.playerY[-2] ),
    .A1(\rbzero.debug_overlay.playerX[-2] ),
    .S(_08138_),
    .X(_09594_));
 sky130_fd_sc_hd__nor2_1 _16504_ (.A(_09593_),
    .B(_09594_),
    .Y(_09595_));
 sky130_fd_sc_hd__and2_1 _16505_ (.A(_09593_),
    .B(_09594_),
    .X(_09596_));
 sky130_fd_sc_hd__nor2_1 _16506_ (.A(_09595_),
    .B(_09596_),
    .Y(_09597_));
 sky130_fd_sc_hd__xor2_1 _16507_ (.A(_09121_),
    .B(_09597_),
    .X(_09598_));
 sky130_fd_sc_hd__xnor2_1 _16508_ (.A(_09477_),
    .B(_09598_),
    .Y(_09599_));
 sky130_fd_sc_hd__or2_1 _16509_ (.A(\rbzero.texu_hot[4] ),
    .B(_08145_),
    .X(_09600_));
 sky130_fd_sc_hd__o211a_1 _16510_ (.A1(_08148_),
    .A2(_09599_),
    .B1(_09600_),
    .C1(_08085_),
    .X(_00470_));
 sky130_fd_sc_hd__o21ba_1 _16511_ (.A1(_09477_),
    .A2(_09595_),
    .B1_N(_09596_),
    .X(_09601_));
 sky130_fd_sc_hd__o21a_1 _16512_ (.A1(_09479_),
    .A2(_09592_),
    .B1(_09590_),
    .X(_09602_));
 sky130_fd_sc_hd__or2b_1 _16513_ (.A(_09513_),
    .B_N(_09484_),
    .X(_09603_));
 sky130_fd_sc_hd__or2b_1 _16514_ (.A(_09487_),
    .B_N(_09494_),
    .X(_09604_));
 sky130_fd_sc_hd__a21oi_1 _16515_ (.A1(_09511_),
    .A2(_09603_),
    .B1(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__and3_1 _16516_ (.A(_09604_),
    .B(_09511_),
    .C(_09603_),
    .X(_09606_));
 sky130_fd_sc_hd__nor2_1 _16517_ (.A(_09605_),
    .B(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__nand2_1 _16518_ (.A(\rbzero.wall_tracer.visualWallDist[10] ),
    .B(_08475_),
    .Y(_09608_));
 sky130_fd_sc_hd__or2_2 _16519_ (.A(_08170_),
    .B(_09608_),
    .X(_09609_));
 sky130_fd_sc_hd__xnor2_1 _16520_ (.A(_09607_),
    .B(_09609_),
    .Y(_09610_));
 sky130_fd_sc_hd__a21o_1 _16521_ (.A1(_09495_),
    .A2(_09509_),
    .B1(_09507_),
    .X(_09611_));
 sky130_fd_sc_hd__or2b_1 _16522_ (.A(_09539_),
    .B_N(_09518_),
    .X(_09612_));
 sky130_fd_sc_hd__or2b_1 _16523_ (.A(_09540_),
    .B_N(_09515_),
    .X(_09613_));
 sky130_fd_sc_hd__nor2_1 _16524_ (.A(_09008_),
    .B(_09363_),
    .Y(_09614_));
 sky130_fd_sc_hd__nor2_1 _16525_ (.A(_09005_),
    .B(_09242_),
    .Y(_09615_));
 sky130_fd_sc_hd__o22a_1 _16526_ (.A1(_09005_),
    .A2(_09252_),
    .B1(_09243_),
    .B2(_08952_),
    .X(_09616_));
 sky130_fd_sc_hd__a21oi_1 _16527_ (.A1(_09498_),
    .A2(_09615_),
    .B1(_09616_),
    .Y(_09617_));
 sky130_fd_sc_hd__xnor2_1 _16528_ (.A(_09614_),
    .B(_09617_),
    .Y(_09618_));
 sky130_fd_sc_hd__a21oi_1 _16529_ (.A1(_09365_),
    .A2(_09614_),
    .B1(_09492_),
    .Y(_09619_));
 sky130_fd_sc_hd__xor2_1 _16530_ (.A(_09618_),
    .B(_09619_),
    .X(_09620_));
 sky130_fd_sc_hd__buf_4 _16531_ (.A(_09491_),
    .X(_09621_));
 sky130_fd_sc_hd__nor2_1 _16532_ (.A(_08304_),
    .B(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__xor2_1 _16533_ (.A(_09620_),
    .B(_09622_),
    .X(_09623_));
 sky130_fd_sc_hd__nand2_1 _16534_ (.A(_09371_),
    .B(_09499_),
    .Y(_09624_));
 sky130_fd_sc_hd__a21bo_1 _16535_ (.A1(_09498_),
    .A2(_09501_),
    .B1_N(_09624_),
    .X(_09625_));
 sky130_fd_sc_hd__a21bo_1 _16536_ (.A1(_09521_),
    .A2(_09526_),
    .B1_N(_09523_),
    .X(_09626_));
 sky130_fd_sc_hd__o22a_1 _16537_ (.A1(_09520_),
    .A2(_08541_),
    .B1(_08618_),
    .B2(_09525_),
    .X(_09627_));
 sky130_fd_sc_hd__or2_1 _16538_ (.A(_08734_),
    .B(_08617_),
    .X(_09628_));
 sky130_fd_sc_hd__or3_1 _16539_ (.A(_08731_),
    .B(_08541_),
    .C(_09628_),
    .X(_09629_));
 sky130_fd_sc_hd__and2b_1 _16540_ (.A_N(_09627_),
    .B(_09629_),
    .X(_09630_));
 sky130_fd_sc_hd__xor2_1 _16541_ (.A(_09499_),
    .B(_09630_),
    .X(_09631_));
 sky130_fd_sc_hd__xor2_1 _16542_ (.A(_09626_),
    .B(_09631_),
    .X(_09632_));
 sky130_fd_sc_hd__xnor2_1 _16543_ (.A(_09625_),
    .B(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__a21oi_1 _16544_ (.A1(_09497_),
    .A2(_09505_),
    .B1(_09503_),
    .Y(_09634_));
 sky130_fd_sc_hd__nor2_1 _16545_ (.A(_09633_),
    .B(_09634_),
    .Y(_09635_));
 sky130_fd_sc_hd__nand2_1 _16546_ (.A(_09633_),
    .B(_09634_),
    .Y(_09636_));
 sky130_fd_sc_hd__and2b_1 _16547_ (.A_N(_09635_),
    .B(_09636_),
    .X(_09637_));
 sky130_fd_sc_hd__xnor2_1 _16548_ (.A(_09623_),
    .B(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__a21o_1 _16549_ (.A1(_09612_),
    .A2(_09613_),
    .B1(_09638_),
    .X(_09639_));
 sky130_fd_sc_hd__nand3_1 _16550_ (.A(_09612_),
    .B(_09613_),
    .C(_09638_),
    .Y(_09640_));
 sky130_fd_sc_hd__nand2_1 _16551_ (.A(_09639_),
    .B(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__xnor2_1 _16552_ (.A(_09611_),
    .B(_09641_),
    .Y(_09642_));
 sky130_fd_sc_hd__a21o_1 _16553_ (.A1(_09527_),
    .A2(_09537_),
    .B1(_09536_),
    .X(_09643_));
 sky130_fd_sc_hd__nand2_1 _16554_ (.A(_09546_),
    .B(_09552_),
    .Y(_09644_));
 sky130_fd_sc_hd__a21bo_1 _16555_ (.A1(_09544_),
    .A2(_09553_),
    .B1_N(_09644_),
    .X(_09645_));
 sky130_fd_sc_hd__or4_1 _16556_ (.A(_08152_),
    .B(_08535_),
    .C(_08409_),
    .D(_08382_),
    .X(_09646_));
 sky130_fd_sc_hd__clkbuf_4 _16557_ (.A(_08382_),
    .X(_09647_));
 sky130_fd_sc_hd__o22ai_1 _16558_ (.A1(_08535_),
    .A2(_08409_),
    .B1(_09647_),
    .B2(_08152_),
    .Y(_09648_));
 sky130_fd_sc_hd__nand2_1 _16559_ (.A(_09646_),
    .B(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__xor2_1 _16560_ (.A(_09522_),
    .B(_09649_),
    .X(_09650_));
 sky130_fd_sc_hd__or2_1 _16561_ (.A(_08813_),
    .B(_09037_),
    .X(_09651_));
 sky130_fd_sc_hd__o22ai_1 _16562_ (.A1(_08813_),
    .A2(_09176_),
    .B1(_09037_),
    .B2(_09406_),
    .Y(_09652_));
 sky130_fd_sc_hd__o31a_1 _16563_ (.A1(_09406_),
    .A2(_09176_),
    .A3(_09651_),
    .B1(_09652_),
    .X(_09653_));
 sky130_fd_sc_hd__xnor2_1 _16564_ (.A(_09529_),
    .B(_09653_),
    .Y(_09654_));
 sky130_fd_sc_hd__a22oi_2 _16565_ (.A1(_09393_),
    .A2(_09529_),
    .B1(_09531_),
    .B2(_09532_),
    .Y(_09655_));
 sky130_fd_sc_hd__nor2_1 _16566_ (.A(_09654_),
    .B(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__nand2_1 _16567_ (.A(_09654_),
    .B(_09655_),
    .Y(_09657_));
 sky130_fd_sc_hd__and2b_1 _16568_ (.A_N(_09656_),
    .B(_09657_),
    .X(_09658_));
 sky130_fd_sc_hd__xnor2_1 _16569_ (.A(_09650_),
    .B(_09658_),
    .Y(_09659_));
 sky130_fd_sc_hd__xor2_1 _16570_ (.A(_09645_),
    .B(_09659_),
    .X(_09660_));
 sky130_fd_sc_hd__xnor2_1 _16571_ (.A(_09643_),
    .B(_09660_),
    .Y(_09661_));
 sky130_fd_sc_hd__clkbuf_4 _16572_ (.A(_09044_),
    .X(_09662_));
 sky130_fd_sc_hd__a21oi_1 _16573_ (.A1(_09662_),
    .A2(_09046_),
    .B1(_08816_),
    .Y(_09663_));
 sky130_fd_sc_hd__a21bo_1 _16574_ (.A1(_09410_),
    .A2(_09663_),
    .B1_N(_09550_),
    .X(_09664_));
 sky130_fd_sc_hd__or3_1 _16575_ (.A(_09167_),
    .B(_09186_),
    .C(_09556_),
    .X(_09665_));
 sky130_fd_sc_hd__a21bo_1 _16576_ (.A1(_09545_),
    .A2(_09555_),
    .B1_N(_09665_),
    .X(_09666_));
 sky130_fd_sc_hd__a21oi_2 _16577_ (.A1(_09315_),
    .A2(_09306_),
    .B1(_08369_),
    .Y(_09667_));
 sky130_fd_sc_hd__and2_1 _16578_ (.A(_09053_),
    .B(_09306_),
    .X(_09668_));
 sky130_fd_sc_hd__buf_2 _16579_ (.A(_09668_),
    .X(_09669_));
 sky130_fd_sc_hd__clkbuf_4 _16580_ (.A(_08466_),
    .X(_09670_));
 sky130_fd_sc_hd__a21oi_1 _16581_ (.A1(_09670_),
    .A2(_09184_),
    .B1(_08889_),
    .Y(_09671_));
 sky130_fd_sc_hd__o21ba_1 _16582_ (.A1(_08434_),
    .A2(_09669_),
    .B1_N(_09671_),
    .X(_09672_));
 sky130_fd_sc_hd__a21oi_1 _16583_ (.A1(_09557_),
    .A2(_09667_),
    .B1(_09672_),
    .Y(_09673_));
 sky130_fd_sc_hd__xor2_1 _16584_ (.A(_09663_),
    .B(_09673_),
    .X(_09674_));
 sky130_fd_sc_hd__xor2_1 _16585_ (.A(_09666_),
    .B(_09674_),
    .X(_09675_));
 sky130_fd_sc_hd__xor2_1 _16586_ (.A(_09664_),
    .B(_09675_),
    .X(_09676_));
 sky130_fd_sc_hd__buf_2 _16587_ (.A(_09422_),
    .X(_09677_));
 sky130_fd_sc_hd__nor2_1 _16588_ (.A(_08910_),
    .B(_09677_),
    .Y(_09678_));
 sky130_fd_sc_hd__or2_1 _16589_ (.A(_08950_),
    .B(_09559_),
    .X(_09679_));
 sky130_fd_sc_hd__mux2_2 _16590_ (.A0(\rbzero.wall_tracer.stepDistX[8] ),
    .A1(_09426_),
    .S(_06263_),
    .X(_09680_));
 sky130_fd_sc_hd__nand2b_2 _16591_ (.A_N(_08431_),
    .B(_09680_),
    .Y(_09681_));
 sky130_fd_sc_hd__a2bb2o_1 _16592_ (.A1_N(_08431_),
    .A2_N(_09559_),
    .B1(_09680_),
    .B2(_08733_),
    .X(_09682_));
 sky130_fd_sc_hd__o21a_1 _16593_ (.A1(_09679_),
    .A2(_09681_),
    .B1(_09682_),
    .X(_09683_));
 sky130_fd_sc_hd__xor2_1 _16594_ (.A(_09678_),
    .B(_09683_),
    .X(_09684_));
 sky130_fd_sc_hd__nand2_1 _16595_ (.A(\rbzero.wall_tracer.stepDistY[9] ),
    .B(_08405_),
    .Y(_09685_));
 sky130_fd_sc_hd__a21oi_2 _16596_ (.A1(_09685_),
    .A2(_09566_),
    .B1(_08458_),
    .Y(_09686_));
 sky130_fd_sc_hd__nor2_2 _16597_ (.A(_06433_),
    .B(_08338_),
    .Y(_09687_));
 sky130_fd_sc_hd__or4_1 _16598_ (.A(_08027_),
    .B(_08029_),
    .C(_08031_),
    .D(_09563_),
    .X(_09688_));
 sky130_fd_sc_hd__a21o_1 _16599_ (.A1(_08148_),
    .A2(_09688_),
    .B1(_08454_),
    .X(_09689_));
 sky130_fd_sc_hd__or3_1 _16600_ (.A(_08039_),
    .B(_08338_),
    .C(_09689_),
    .X(_09690_));
 sky130_fd_sc_hd__buf_2 _16601_ (.A(_09690_),
    .X(_09691_));
 sky130_fd_sc_hd__mux2_1 _16602_ (.A0(_06433_),
    .A1(_09687_),
    .S(_09691_),
    .X(_09692_));
 sky130_fd_sc_hd__xnor2_1 _16603_ (.A(_09686_),
    .B(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__nor2_1 _16604_ (.A(_09562_),
    .B(_09567_),
    .Y(_09694_));
 sky130_fd_sc_hd__a21oi_1 _16605_ (.A1(_09561_),
    .A2(_09568_),
    .B1(_09694_),
    .Y(_09695_));
 sky130_fd_sc_hd__xor2_1 _16606_ (.A(_09693_),
    .B(_09695_),
    .X(_09696_));
 sky130_fd_sc_hd__xnor2_1 _16607_ (.A(_09684_),
    .B(_09696_),
    .Y(_09697_));
 sky130_fd_sc_hd__and2b_1 _16608_ (.A_N(_09569_),
    .B(_09570_),
    .X(_09698_));
 sky130_fd_sc_hd__a21o_1 _16609_ (.A1(_09558_),
    .A2(_09571_),
    .B1(_09698_),
    .X(_09699_));
 sky130_fd_sc_hd__xnor2_1 _16610_ (.A(_09697_),
    .B(_09699_),
    .Y(_09700_));
 sky130_fd_sc_hd__xnor2_1 _16611_ (.A(_09676_),
    .B(_09700_),
    .Y(_09701_));
 sky130_fd_sc_hd__nor2_1 _16612_ (.A(_09572_),
    .B(_09573_),
    .Y(_09702_));
 sky130_fd_sc_hd__a21o_1 _16613_ (.A1(_09554_),
    .A2(_09574_),
    .B1(_09702_),
    .X(_09703_));
 sky130_fd_sc_hd__xnor2_1 _16614_ (.A(_09701_),
    .B(_09703_),
    .Y(_09704_));
 sky130_fd_sc_hd__xnor2_1 _16615_ (.A(_09661_),
    .B(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__nor2_1 _16616_ (.A(_09575_),
    .B(_09576_),
    .Y(_09706_));
 sky130_fd_sc_hd__a21oi_1 _16617_ (.A1(_09541_),
    .A2(_09577_),
    .B1(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__nor2_1 _16618_ (.A(_09705_),
    .B(_09707_),
    .Y(_09708_));
 sky130_fd_sc_hd__nand2_1 _16619_ (.A(_09705_),
    .B(_09707_),
    .Y(_09709_));
 sky130_fd_sc_hd__and2b_1 _16620_ (.A_N(_09708_),
    .B(_09709_),
    .X(_09710_));
 sky130_fd_sc_hd__xnor2_1 _16621_ (.A(_09642_),
    .B(_09710_),
    .Y(_09711_));
 sky130_fd_sc_hd__a21oi_1 _16622_ (.A1(_09514_),
    .A2(_09581_),
    .B1(_09580_),
    .Y(_09712_));
 sky130_fd_sc_hd__xor2_1 _16623_ (.A(_09711_),
    .B(_09712_),
    .X(_09713_));
 sky130_fd_sc_hd__xnor2_1 _16624_ (.A(_09610_),
    .B(_09713_),
    .Y(_09714_));
 sky130_fd_sc_hd__nor2_1 _16625_ (.A(_09583_),
    .B(_09584_),
    .Y(_09715_));
 sky130_fd_sc_hd__a21oi_1 _16626_ (.A1(_09483_),
    .A2(_09585_),
    .B1(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__nor2_2 _16627_ (.A(_09714_),
    .B(_09716_),
    .Y(_09717_));
 sky130_fd_sc_hd__and2_1 _16628_ (.A(_09714_),
    .B(_09716_),
    .X(_09718_));
 sky130_fd_sc_hd__or2_2 _16629_ (.A(_09717_),
    .B(_09718_),
    .X(_09719_));
 sky130_fd_sc_hd__xor2_4 _16630_ (.A(_09587_),
    .B(_09719_),
    .X(_09720_));
 sky130_fd_sc_hd__xnor2_4 _16631_ (.A(_09602_),
    .B(_09720_),
    .Y(_09721_));
 sky130_fd_sc_hd__mux2_1 _16632_ (.A0(\rbzero.debug_overlay.playerY[-1] ),
    .A1(\rbzero.debug_overlay.playerX[-1] ),
    .S(_08138_),
    .X(_09722_));
 sky130_fd_sc_hd__xnor2_1 _16633_ (.A(_09121_),
    .B(_09722_),
    .Y(_09723_));
 sky130_fd_sc_hd__xnor2_1 _16634_ (.A(_09721_),
    .B(_09723_),
    .Y(_09724_));
 sky130_fd_sc_hd__xnor2_1 _16635_ (.A(_09601_),
    .B(_09724_),
    .Y(_09725_));
 sky130_fd_sc_hd__or2_1 _16636_ (.A(\rbzero.texu_hot[5] ),
    .B(_08145_),
    .X(_09726_));
 sky130_fd_sc_hd__o211a_1 _16637_ (.A1(_08148_),
    .A2(_09725_),
    .B1(_09726_),
    .C1(_04442_),
    .X(_00471_));
 sky130_fd_sc_hd__nor2_1 _16638_ (.A(_04414_),
    .B(_04699_),
    .Y(_09727_));
 sky130_fd_sc_hd__and4_1 _16639_ (.A(_04051_),
    .B(_04637_),
    .C(_05053_),
    .D(_09727_),
    .X(_09728_));
 sky130_fd_sc_hd__clkbuf_4 _16640_ (.A(_09728_),
    .X(_09729_));
 sky130_fd_sc_hd__or2_1 _16641_ (.A(_04408_),
    .B(_09729_),
    .X(_09730_));
 sky130_fd_sc_hd__nor2_1 _16642_ (.A(_03971_),
    .B(_09730_),
    .Y(_00472_));
 sky130_fd_sc_hd__nor2_1 _16643_ (.A(_04408_),
    .B(_09729_),
    .Y(_09731_));
 sky130_fd_sc_hd__clkbuf_4 _16644_ (.A(_09731_),
    .X(_09732_));
 sky130_fd_sc_hd__and3_1 _16645_ (.A(_04447_),
    .B(_04448_),
    .C(_09732_),
    .X(_09733_));
 sky130_fd_sc_hd__clkbuf_1 _16646_ (.A(_09733_),
    .X(_00473_));
 sky130_fd_sc_hd__buf_6 _16647_ (.A(_04408_),
    .X(_09734_));
 sky130_fd_sc_hd__or2_1 _16648_ (.A(_09734_),
    .B(_04636_),
    .X(_09735_));
 sky130_fd_sc_hd__a21oi_1 _16649_ (.A1(_04446_),
    .A2(_04448_),
    .B1(_09735_),
    .Y(_00474_));
 sky130_fd_sc_hd__nor2_1 _16650_ (.A(net63),
    .B(_05061_),
    .Y(_00475_));
 sky130_fd_sc_hd__and3_1 _16651_ (.A(_04638_),
    .B(_05079_),
    .C(_09732_),
    .X(_09736_));
 sky130_fd_sc_hd__clkbuf_1 _16652_ (.A(_09736_),
    .X(_00476_));
 sky130_fd_sc_hd__nor2_1 _16653_ (.A(_05075_),
    .B(_09730_),
    .Y(_00477_));
 sky130_fd_sc_hd__and2_1 _16654_ (.A(_05069_),
    .B(_09732_),
    .X(_09737_));
 sky130_fd_sc_hd__clkbuf_1 _16655_ (.A(_09737_),
    .X(_00478_));
 sky130_fd_sc_hd__and2_1 _16656_ (.A(_05073_),
    .B(_09732_),
    .X(_09738_));
 sky130_fd_sc_hd__clkbuf_1 _16657_ (.A(_09738_),
    .X(_00479_));
 sky130_fd_sc_hd__and4_1 _16658_ (.A(_03975_),
    .B(_04415_),
    .C(_04636_),
    .D(_05283_),
    .X(_09739_));
 sky130_fd_sc_hd__a31o_1 _16659_ (.A1(_04415_),
    .A2(_04636_),
    .A3(_05283_),
    .B1(_03975_),
    .X(_09740_));
 sky130_fd_sc_hd__and3b_1 _16660_ (.A_N(_09739_),
    .B(_09740_),
    .C(_09732_),
    .X(_09741_));
 sky130_fd_sc_hd__clkbuf_1 _16661_ (.A(_09741_),
    .X(_00480_));
 sky130_fd_sc_hd__a21oi_1 _16662_ (.A1(_04420_),
    .A2(_09739_),
    .B1(_09730_),
    .Y(_09742_));
 sky130_fd_sc_hd__o21a_1 _16663_ (.A1(_04420_),
    .A2(_09739_),
    .B1(_09742_),
    .X(_00481_));
 sky130_fd_sc_hd__and3_2 _16664_ (.A(\rbzero.trace_state[0] ),
    .B(_05050_),
    .C(_09729_),
    .X(_09743_));
 sky130_fd_sc_hd__nor2_4 _16665_ (.A(_08134_),
    .B(_09743_),
    .Y(_09744_));
 sky130_fd_sc_hd__clkbuf_4 _16666_ (.A(_09744_),
    .X(_09745_));
 sky130_fd_sc_hd__buf_4 _16667_ (.A(_09745_),
    .X(_09746_));
 sky130_fd_sc_hd__and4_1 _16668_ (.A(_04051_),
    .B(_04637_),
    .C(_05053_),
    .D(_09727_),
    .X(_09747_));
 sky130_fd_sc_hd__and4_1 _16669_ (.A(_04437_),
    .B(_04433_),
    .C(_05050_),
    .D(_09747_),
    .X(_09748_));
 sky130_fd_sc_hd__buf_4 _16670_ (.A(_09748_),
    .X(_09749_));
 sky130_fd_sc_hd__clkbuf_4 _16671_ (.A(_09749_),
    .X(_09750_));
 sky130_fd_sc_hd__a22o_1 _16672_ (.A1(\rbzero.row_render.side ),
    .A2(_09746_),
    .B1(_09750_),
    .B2(_08138_),
    .X(_00482_));
 sky130_fd_sc_hd__a22o_1 _16673_ (.A1(\rbzero.row_render.size[0] ),
    .A2(_09746_),
    .B1(_09750_),
    .B2(_07923_),
    .X(_00483_));
 sky130_fd_sc_hd__a22o_1 _16674_ (.A1(\rbzero.row_render.size[1] ),
    .A2(_09746_),
    .B1(_09750_),
    .B2(_07935_),
    .X(_00484_));
 sky130_fd_sc_hd__a22o_1 _16675_ (.A1(\rbzero.row_render.size[2] ),
    .A2(_09746_),
    .B1(_09750_),
    .B2(_07944_),
    .X(_00485_));
 sky130_fd_sc_hd__a22o_1 _16676_ (.A1(\rbzero.row_render.size[3] ),
    .A2(_09746_),
    .B1(_09750_),
    .B2(_07954_),
    .X(_00486_));
 sky130_fd_sc_hd__a22o_1 _16677_ (.A1(\rbzero.row_render.size[4] ),
    .A2(_09746_),
    .B1(_09750_),
    .B2(_07964_),
    .X(_00487_));
 sky130_fd_sc_hd__a22o_1 _16678_ (.A1(\rbzero.row_render.size[5] ),
    .A2(_09746_),
    .B1(_09750_),
    .B2(_07971_),
    .X(_00488_));
 sky130_fd_sc_hd__a22o_1 _16679_ (.A1(\rbzero.row_render.size[6] ),
    .A2(_09746_),
    .B1(_09750_),
    .B2(_07975_),
    .X(_00489_));
 sky130_fd_sc_hd__clkbuf_8 _16680_ (.A(_09744_),
    .X(_09751_));
 sky130_fd_sc_hd__buf_4 _16681_ (.A(_09751_),
    .X(_09752_));
 sky130_fd_sc_hd__a22o_1 _16682_ (.A1(\rbzero.row_render.size[7] ),
    .A2(_09752_),
    .B1(_09750_),
    .B2(_07982_),
    .X(_00490_));
 sky130_fd_sc_hd__buf_4 _16683_ (.A(_09749_),
    .X(_09753_));
 sky130_fd_sc_hd__buf_4 _16684_ (.A(_09753_),
    .X(_09754_));
 sky130_fd_sc_hd__a22o_1 _16685_ (.A1(\rbzero.row_render.size[8] ),
    .A2(_09752_),
    .B1(_09754_),
    .B2(_07992_),
    .X(_00491_));
 sky130_fd_sc_hd__a22o_1 _16686_ (.A1(\rbzero.row_render.size[9] ),
    .A2(_09752_),
    .B1(_09754_),
    .B2(_07996_),
    .X(_00492_));
 sky130_fd_sc_hd__a22o_1 _16687_ (.A1(\rbzero.row_render.size[10] ),
    .A2(_09752_),
    .B1(_09754_),
    .B2(_08000_),
    .X(_00493_));
 sky130_fd_sc_hd__a22o_1 _16688_ (.A1(\rbzero.row_render.texu[0] ),
    .A2(_09752_),
    .B1(_09754_),
    .B2(\rbzero.texu_hot[0] ),
    .X(_00494_));
 sky130_fd_sc_hd__a22o_1 _16689_ (.A1(\rbzero.row_render.texu[1] ),
    .A2(_09752_),
    .B1(_09754_),
    .B2(\rbzero.texu_hot[1] ),
    .X(_00495_));
 sky130_fd_sc_hd__a22o_1 _16690_ (.A1(\rbzero.row_render.texu[2] ),
    .A2(_09752_),
    .B1(_09754_),
    .B2(\rbzero.texu_hot[2] ),
    .X(_00496_));
 sky130_fd_sc_hd__a22o_1 _16691_ (.A1(\rbzero.row_render.texu[3] ),
    .A2(_09752_),
    .B1(_09754_),
    .B2(\rbzero.texu_hot[3] ),
    .X(_00497_));
 sky130_fd_sc_hd__a22o_1 _16692_ (.A1(\rbzero.row_render.texu[4] ),
    .A2(_09752_),
    .B1(_09754_),
    .B2(\rbzero.texu_hot[4] ),
    .X(_00498_));
 sky130_fd_sc_hd__a22o_1 _16693_ (.A1(\rbzero.traced_texa[-11] ),
    .A2(_09752_),
    .B1(_09754_),
    .B2(\rbzero.wall_tracer.visualWallDist[-11] ),
    .X(_00499_));
 sky130_fd_sc_hd__clkbuf_4 _16694_ (.A(_09751_),
    .X(_09755_));
 sky130_fd_sc_hd__a22o_1 _16695_ (.A1(\rbzero.traced_texa[-10] ),
    .A2(_09755_),
    .B1(_09754_),
    .B2(\rbzero.wall_tracer.visualWallDist[-10] ),
    .X(_00500_));
 sky130_fd_sc_hd__clkbuf_4 _16696_ (.A(_09753_),
    .X(_09756_));
 sky130_fd_sc_hd__a22o_1 _16697_ (.A1(\rbzero.traced_texa[-9] ),
    .A2(_09755_),
    .B1(_09756_),
    .B2(\rbzero.wall_tracer.visualWallDist[-9] ),
    .X(_00501_));
 sky130_fd_sc_hd__a22o_1 _16698_ (.A1(\rbzero.traced_texa[-8] ),
    .A2(_09755_),
    .B1(_09756_),
    .B2(\rbzero.wall_tracer.visualWallDist[-8] ),
    .X(_00502_));
 sky130_fd_sc_hd__a22o_1 _16699_ (.A1(\rbzero.traced_texa[-7] ),
    .A2(_09755_),
    .B1(_09756_),
    .B2(\rbzero.wall_tracer.visualWallDist[-7] ),
    .X(_00503_));
 sky130_fd_sc_hd__a22o_1 _16700_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(_09755_),
    .B1(_09756_),
    .B2(\rbzero.wall_tracer.visualWallDist[-6] ),
    .X(_00504_));
 sky130_fd_sc_hd__a22o_1 _16701_ (.A1(\rbzero.traced_texa[-5] ),
    .A2(_09755_),
    .B1(_09756_),
    .B2(\rbzero.wall_tracer.visualWallDist[-5] ),
    .X(_00505_));
 sky130_fd_sc_hd__a22o_1 _16702_ (.A1(\rbzero.traced_texa[-4] ),
    .A2(_09755_),
    .B1(_09756_),
    .B2(\rbzero.wall_tracer.visualWallDist[-4] ),
    .X(_00506_));
 sky130_fd_sc_hd__a22o_1 _16703_ (.A1(\rbzero.traced_texa[-3] ),
    .A2(_09755_),
    .B1(_09756_),
    .B2(\rbzero.wall_tracer.visualWallDist[-3] ),
    .X(_00507_));
 sky130_fd_sc_hd__a22o_1 _16704_ (.A1(\rbzero.traced_texa[-2] ),
    .A2(_09755_),
    .B1(_09756_),
    .B2(\rbzero.wall_tracer.visualWallDist[-2] ),
    .X(_00508_));
 sky130_fd_sc_hd__a22o_1 _16705_ (.A1(\rbzero.traced_texa[-1] ),
    .A2(_09755_),
    .B1(_09756_),
    .B2(\rbzero.wall_tracer.visualWallDist[-1] ),
    .X(_00509_));
 sky130_fd_sc_hd__clkbuf_4 _16706_ (.A(_09751_),
    .X(_09757_));
 sky130_fd_sc_hd__a22o_1 _16707_ (.A1(\rbzero.traced_texa[0] ),
    .A2(_09757_),
    .B1(_09756_),
    .B2(\rbzero.wall_tracer.visualWallDist[0] ),
    .X(_00510_));
 sky130_fd_sc_hd__buf_2 _16708_ (.A(_09749_),
    .X(_09758_));
 sky130_fd_sc_hd__a22o_1 _16709_ (.A1(\rbzero.traced_texa[1] ),
    .A2(_09757_),
    .B1(_09758_),
    .B2(\rbzero.wall_tracer.visualWallDist[1] ),
    .X(_00511_));
 sky130_fd_sc_hd__a22o_1 _16710_ (.A1(\rbzero.traced_texa[2] ),
    .A2(_09757_),
    .B1(_09758_),
    .B2(\rbzero.wall_tracer.visualWallDist[2] ),
    .X(_00512_));
 sky130_fd_sc_hd__a22o_1 _16711_ (.A1(\rbzero.traced_texa[3] ),
    .A2(_09757_),
    .B1(_09758_),
    .B2(\rbzero.wall_tracer.visualWallDist[3] ),
    .X(_00513_));
 sky130_fd_sc_hd__a22o_1 _16712_ (.A1(\rbzero.traced_texa[4] ),
    .A2(_09757_),
    .B1(_09758_),
    .B2(\rbzero.wall_tracer.visualWallDist[4] ),
    .X(_00514_));
 sky130_fd_sc_hd__a22o_1 _16713_ (.A1(\rbzero.traced_texa[5] ),
    .A2(_09757_),
    .B1(_09758_),
    .B2(\rbzero.wall_tracer.visualWallDist[5] ),
    .X(_00515_));
 sky130_fd_sc_hd__a22o_1 _16714_ (.A1(\rbzero.traced_texa[6] ),
    .A2(_09757_),
    .B1(_09758_),
    .B2(\rbzero.wall_tracer.visualWallDist[6] ),
    .X(_00516_));
 sky130_fd_sc_hd__a22o_1 _16715_ (.A1(\rbzero.traced_texa[7] ),
    .A2(_09757_),
    .B1(_09758_),
    .B2(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_00517_));
 sky130_fd_sc_hd__a22o_1 _16716_ (.A1(\rbzero.traced_texa[8] ),
    .A2(_09757_),
    .B1(_09758_),
    .B2(\rbzero.wall_tracer.visualWallDist[8] ),
    .X(_00518_));
 sky130_fd_sc_hd__a22o_1 _16717_ (.A1(\rbzero.traced_texa[9] ),
    .A2(_09757_),
    .B1(_09758_),
    .B2(\rbzero.wall_tracer.visualWallDist[9] ),
    .X(_00519_));
 sky130_fd_sc_hd__buf_2 _16718_ (.A(_09751_),
    .X(_09759_));
 sky130_fd_sc_hd__a22o_1 _16719_ (.A1(\rbzero.traced_texa[10] ),
    .A2(_09759_),
    .B1(_09758_),
    .B2(\rbzero.wall_tracer.visualWallDist[10] ),
    .X(_00520_));
 sky130_fd_sc_hd__nand4_4 _16720_ (.A(_04437_),
    .B(_04433_),
    .C(_05050_),
    .D(_09729_),
    .Y(_09760_));
 sky130_fd_sc_hd__mux2_1 _16721_ (.A0(\rbzero.wall_hot[0] ),
    .A1(\rbzero.row_render.wall[0] ),
    .S(_09760_),
    .X(_09761_));
 sky130_fd_sc_hd__clkbuf_1 _16722_ (.A(_09761_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _16723_ (.A0(\rbzero.wall_hot[1] ),
    .A1(\rbzero.row_render.wall[1] ),
    .S(_09760_),
    .X(_09762_));
 sky130_fd_sc_hd__clkbuf_1 _16724_ (.A(_09762_),
    .X(_00522_));
 sky130_fd_sc_hd__o21a_1 _16725_ (.A1(\rbzero.map_rom.i_col[4] ),
    .A2(\rbzero.wall_tracer.mapX[5] ),
    .B1(_09118_),
    .X(_09763_));
 sky130_fd_sc_hd__xnor2_1 _16726_ (.A(_06126_),
    .B(_09118_),
    .Y(_09764_));
 sky130_fd_sc_hd__and2_1 _16727_ (.A(\rbzero.map_rom.f1 ),
    .B(_09118_),
    .X(_09765_));
 sky130_fd_sc_hd__xnor2_1 _16728_ (.A(_06117_),
    .B(_08218_),
    .Y(_09766_));
 sky130_fd_sc_hd__and2_1 _16729_ (.A(\rbzero.map_rom.f4 ),
    .B(_09766_),
    .X(_09767_));
 sky130_fd_sc_hd__a21o_1 _16730_ (.A1(_06113_),
    .A2(_09118_),
    .B1(_09767_),
    .X(_09768_));
 sky130_fd_sc_hd__and2_1 _16731_ (.A(\rbzero.map_rom.f2 ),
    .B(_08218_),
    .X(_09769_));
 sky130_fd_sc_hd__nor2_1 _16732_ (.A(\rbzero.map_rom.f2 ),
    .B(_08218_),
    .Y(_09770_));
 sky130_fd_sc_hd__nor2_1 _16733_ (.A(_09769_),
    .B(_09770_),
    .Y(_09771_));
 sky130_fd_sc_hd__a21o_1 _16734_ (.A1(_09768_),
    .A2(_09771_),
    .B1(_09769_),
    .X(_09772_));
 sky130_fd_sc_hd__or2_1 _16735_ (.A(\rbzero.map_rom.f1 ),
    .B(_09118_),
    .X(_09773_));
 sky130_fd_sc_hd__o21ai_1 _16736_ (.A1(_09765_),
    .A2(_09772_),
    .B1(_09773_),
    .Y(_09774_));
 sky130_fd_sc_hd__xnor2_1 _16737_ (.A(_06129_),
    .B(_09118_),
    .Y(_09775_));
 sky130_fd_sc_hd__and2b_1 _16738_ (.A_N(_09774_),
    .B(_09775_),
    .X(_09776_));
 sky130_fd_sc_hd__and2_1 _16739_ (.A(_09764_),
    .B(_09776_),
    .X(_09777_));
 sky130_fd_sc_hd__xor2_1 _16740_ (.A(\rbzero.wall_tracer.mapX[6] ),
    .B(_09118_),
    .X(_09778_));
 sky130_fd_sc_hd__o21ai_1 _16741_ (.A1(_09763_),
    .A2(_09777_),
    .B1(_09778_),
    .Y(_09779_));
 sky130_fd_sc_hd__or3_1 _16742_ (.A(_09778_),
    .B(_09763_),
    .C(_09777_),
    .X(_09780_));
 sky130_fd_sc_hd__a21o_1 _16743_ (.A1(_06217_),
    .A2(_06257_),
    .B1(_06161_),
    .X(_09781_));
 sky130_fd_sc_hd__and2_4 _16744_ (.A(_06264_),
    .B(_09781_),
    .X(_09782_));
 sky130_fd_sc_hd__inv_2 _16745_ (.A(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__nor2_2 _16746_ (.A(_06105_),
    .B(_09783_),
    .Y(_09784_));
 sky130_fd_sc_hd__buf_6 _16747_ (.A(_09783_),
    .X(_09785_));
 sky130_fd_sc_hd__a32o_1 _16748_ (.A1(_09779_),
    .A2(_09780_),
    .A3(_09784_),
    .B1(_09785_),
    .B2(\rbzero.wall_tracer.mapX[6] ),
    .X(_00523_));
 sky130_fd_sc_hd__clkbuf_4 _16749_ (.A(_09783_),
    .X(_09786_));
 sky130_fd_sc_hd__xor2_1 _16750_ (.A(\rbzero.wall_tracer.mapX[7] ),
    .B(_09118_),
    .X(_09787_));
 sky130_fd_sc_hd__a21boi_1 _16751_ (.A1(\rbzero.wall_tracer.mapX[6] ),
    .A2(_09119_),
    .B1_N(_09779_),
    .Y(_09788_));
 sky130_fd_sc_hd__xnor2_1 _16752_ (.A(_09787_),
    .B(_09788_),
    .Y(_09789_));
 sky130_fd_sc_hd__a22o_1 _16753_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(_09786_),
    .B1(_09784_),
    .B2(_09789_),
    .X(_00524_));
 sky130_fd_sc_hd__xor2_1 _16754_ (.A(\rbzero.wall_tracer.mapX[8] ),
    .B(_09119_),
    .X(_09790_));
 sky130_fd_sc_hd__and3_1 _16755_ (.A(_09778_),
    .B(_09777_),
    .C(_09787_),
    .X(_09791_));
 sky130_fd_sc_hd__o21a_1 _16756_ (.A1(\rbzero.wall_tracer.mapX[7] ),
    .A2(\rbzero.wall_tracer.mapX[6] ),
    .B1(_09118_),
    .X(_09792_));
 sky130_fd_sc_hd__or3_1 _16757_ (.A(_09763_),
    .B(_09791_),
    .C(_09792_),
    .X(_09793_));
 sky130_fd_sc_hd__xor2_1 _16758_ (.A(_09790_),
    .B(_09793_),
    .X(_09794_));
 sky130_fd_sc_hd__a22o_1 _16759_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_09786_),
    .B1(_09784_),
    .B2(_09794_),
    .X(_00525_));
 sky130_fd_sc_hd__a22o_1 _16760_ (.A1(\rbzero.wall_tracer.mapX[8] ),
    .A2(_09119_),
    .B1(_09790_),
    .B2(_09793_),
    .X(_09795_));
 sky130_fd_sc_hd__xnor2_1 _16761_ (.A(\rbzero.wall_tracer.mapX[9] ),
    .B(_09119_),
    .Y(_09796_));
 sky130_fd_sc_hd__xnor2_1 _16762_ (.A(_09795_),
    .B(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__a22o_1 _16763_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09786_),
    .B1(_09784_),
    .B2(_09797_),
    .X(_00526_));
 sky130_fd_sc_hd__o21a_1 _16764_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09119_),
    .B1(_09795_),
    .X(_09798_));
 sky130_fd_sc_hd__a21oi_1 _16765_ (.A1(\rbzero.wall_tracer.mapX[9] ),
    .A2(_09119_),
    .B1(_09798_),
    .Y(_09799_));
 sky130_fd_sc_hd__xnor2_1 _16766_ (.A(\rbzero.wall_tracer.mapX[10] ),
    .B(_09799_),
    .Y(_09800_));
 sky130_fd_sc_hd__nand2_1 _16767_ (.A(_09119_),
    .B(_09800_),
    .Y(_09801_));
 sky130_fd_sc_hd__or2_1 _16768_ (.A(_09119_),
    .B(_09800_),
    .X(_09802_));
 sky130_fd_sc_hd__a32o_1 _16769_ (.A1(_09784_),
    .A2(_09801_),
    .A3(_09802_),
    .B1(_09785_),
    .B2(\rbzero.wall_tracer.mapX[10] ),
    .X(_00527_));
 sky130_fd_sc_hd__a21oi_1 _16770_ (.A1(_08942_),
    .A2(_08988_),
    .B1(_08123_),
    .Y(_09803_));
 sky130_fd_sc_hd__o21ai_1 _16771_ (.A1(_08942_),
    .A2(_08988_),
    .B1(_09803_),
    .Y(_09804_));
 sky130_fd_sc_hd__o21ai_1 _16772_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_08123_),
    .Y(_09805_));
 sky130_fd_sc_hd__a21o_1 _16773_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09805_),
    .X(_09806_));
 sky130_fd_sc_hd__and3_1 _16774_ (.A(_09782_),
    .B(_09804_),
    .C(_09806_),
    .X(_09807_));
 sky130_fd_sc_hd__a21oi_1 _16775_ (.A1(_06189_),
    .A2(_09786_),
    .B1(_09807_),
    .Y(_00528_));
 sky130_fd_sc_hd__or2_1 _16776_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .X(_09808_));
 sky130_fd_sc_hd__nand2_1 _16777_ (.A(\rbzero.wall_tracer.trackDistX[-10] ),
    .B(\rbzero.wall_tracer.stepDistX[-10] ),
    .Y(_09809_));
 sky130_fd_sc_hd__and4_1 _16778_ (.A(\rbzero.wall_tracer.trackDistX[-11] ),
    .B(\rbzero.wall_tracer.stepDistX[-11] ),
    .C(_09808_),
    .D(_09809_),
    .X(_09810_));
 sky130_fd_sc_hd__a22oi_1 _16779_ (.A1(\rbzero.wall_tracer.trackDistX[-11] ),
    .A2(\rbzero.wall_tracer.stepDistX[-11] ),
    .B1(_09808_),
    .B2(_09809_),
    .Y(_09811_));
 sky130_fd_sc_hd__buf_4 _16780_ (.A(_09782_),
    .X(_09812_));
 sky130_fd_sc_hd__and2_1 _16781_ (.A(_08905_),
    .B(_08990_),
    .X(_09813_));
 sky130_fd_sc_hd__nor2_1 _16782_ (.A(_08905_),
    .B(_08990_),
    .Y(_09814_));
 sky130_fd_sc_hd__or3_1 _16783_ (.A(_08123_),
    .B(_09813_),
    .C(_09814_),
    .X(_09815_));
 sky130_fd_sc_hd__o311a_1 _16784_ (.A1(_06105_),
    .A2(_09810_),
    .A3(_09811_),
    .B1(_09812_),
    .C1(_09815_),
    .X(_09816_));
 sky130_fd_sc_hd__a21oi_1 _16785_ (.A1(_06188_),
    .A2(_09786_),
    .B1(_09816_),
    .Y(_00529_));
 sky130_fd_sc_hd__a21o_1 _16786_ (.A1(\rbzero.wall_tracer.trackDistX[-10] ),
    .A2(\rbzero.wall_tracer.stepDistX[-10] ),
    .B1(_09810_),
    .X(_09817_));
 sky130_fd_sc_hd__or2_1 _16787_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .X(_09818_));
 sky130_fd_sc_hd__nand2_1 _16788_ (.A(\rbzero.wall_tracer.trackDistX[-9] ),
    .B(\rbzero.wall_tracer.stepDistX[-9] ),
    .Y(_09819_));
 sky130_fd_sc_hd__and3_1 _16789_ (.A(_09817_),
    .B(_09818_),
    .C(_09819_),
    .X(_09820_));
 sky130_fd_sc_hd__a21oi_1 _16790_ (.A1(_09818_),
    .A2(_09819_),
    .B1(_09817_),
    .Y(_09821_));
 sky130_fd_sc_hd__clkbuf_4 _16791_ (.A(_06103_),
    .X(_09822_));
 sky130_fd_sc_hd__nand2_1 _16792_ (.A(_09822_),
    .B(_09108_),
    .Y(_09823_));
 sky130_fd_sc_hd__o311a_1 _16793_ (.A1(_06105_),
    .A2(_09820_),
    .A3(_09821_),
    .B1(_09812_),
    .C1(_09823_),
    .X(_09824_));
 sky130_fd_sc_hd__a21oi_1 _16794_ (.A1(_06187_),
    .A2(_09786_),
    .B1(_09824_),
    .Y(_00530_));
 sky130_fd_sc_hd__or2_1 _16795_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .X(_09825_));
 sky130_fd_sc_hd__nand2_1 _16796_ (.A(\rbzero.wall_tracer.trackDistX[-8] ),
    .B(\rbzero.wall_tracer.stepDistX[-8] ),
    .Y(_09826_));
 sky130_fd_sc_hd__a21bo_1 _16797_ (.A1(_09817_),
    .A2(_09818_),
    .B1_N(_09819_),
    .X(_09827_));
 sky130_fd_sc_hd__and3_1 _16798_ (.A(_09825_),
    .B(_09826_),
    .C(_09827_),
    .X(_09828_));
 sky130_fd_sc_hd__a21oi_1 _16799_ (.A1(_09825_),
    .A2(_09826_),
    .B1(_09827_),
    .Y(_09829_));
 sky130_fd_sc_hd__nand2_1 _16800_ (.A(_09822_),
    .B(_09111_),
    .Y(_09830_));
 sky130_fd_sc_hd__o311a_1 _16801_ (.A1(_06105_),
    .A2(_09828_),
    .A3(_09829_),
    .B1(_09812_),
    .C1(_09830_),
    .X(_09831_));
 sky130_fd_sc_hd__a21oi_1 _16802_ (.A1(_06186_),
    .A2(_09786_),
    .B1(_09831_),
    .Y(_00531_));
 sky130_fd_sc_hd__nor2_1 _16803_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_09832_));
 sky130_fd_sc_hd__nand2_1 _16804_ (.A(\rbzero.wall_tracer.trackDistX[-7] ),
    .B(\rbzero.wall_tracer.stepDistX[-7] ),
    .Y(_09833_));
 sky130_fd_sc_hd__or2b_1 _16805_ (.A(_09832_),
    .B_N(_09833_),
    .X(_09834_));
 sky130_fd_sc_hd__a21boi_1 _16806_ (.A1(_09825_),
    .A2(_09827_),
    .B1_N(_09826_),
    .Y(_09835_));
 sky130_fd_sc_hd__xnor2_1 _16807_ (.A(_09834_),
    .B(_09835_),
    .Y(_09836_));
 sky130_fd_sc_hd__nand2_1 _16808_ (.A(_09822_),
    .B(_09105_),
    .Y(_09837_));
 sky130_fd_sc_hd__o211a_1 _16809_ (.A1(_06105_),
    .A2(_09836_),
    .B1(_09837_),
    .C1(_09812_),
    .X(_09838_));
 sky130_fd_sc_hd__a21oi_1 _16810_ (.A1(_06185_),
    .A2(_09786_),
    .B1(_09838_),
    .Y(_00532_));
 sky130_fd_sc_hd__or2_1 _16811_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .X(_09839_));
 sky130_fd_sc_hd__nand2_1 _16812_ (.A(\rbzero.wall_tracer.trackDistX[-6] ),
    .B(\rbzero.wall_tracer.stepDistX[-6] ),
    .Y(_09840_));
 sky130_fd_sc_hd__o21ai_1 _16813_ (.A1(_09832_),
    .A2(_09835_),
    .B1(_09833_),
    .Y(_09841_));
 sky130_fd_sc_hd__a21oi_1 _16814_ (.A1(_09839_),
    .A2(_09840_),
    .B1(_09841_),
    .Y(_09842_));
 sky130_fd_sc_hd__a31o_1 _16815_ (.A1(_09839_),
    .A2(_09840_),
    .A3(_09841_),
    .B1(_06104_),
    .X(_09843_));
 sky130_fd_sc_hd__buf_6 _16816_ (.A(_09782_),
    .X(_09844_));
 sky130_fd_sc_hd__nand2_1 _16817_ (.A(_09822_),
    .B(_09101_),
    .Y(_09845_));
 sky130_fd_sc_hd__o211a_1 _16818_ (.A1(_09842_),
    .A2(_09843_),
    .B1(_09844_),
    .C1(_09845_),
    .X(_09846_));
 sky130_fd_sc_hd__a21oi_1 _16819_ (.A1(_06184_),
    .A2(_09786_),
    .B1(_09846_),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2_1 _16820_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_09847_));
 sky130_fd_sc_hd__nand2_1 _16821_ (.A(\rbzero.wall_tracer.trackDistX[-5] ),
    .B(\rbzero.wall_tracer.stepDistX[-5] ),
    .Y(_09848_));
 sky130_fd_sc_hd__or2b_1 _16822_ (.A(_09847_),
    .B_N(_09848_),
    .X(_09849_));
 sky130_fd_sc_hd__a21boi_1 _16823_ (.A1(_09839_),
    .A2(_09841_),
    .B1_N(_09840_),
    .Y(_09850_));
 sky130_fd_sc_hd__xnor2_1 _16824_ (.A(_09849_),
    .B(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__nand2_1 _16825_ (.A(_06104_),
    .B(_09227_),
    .Y(_09852_));
 sky130_fd_sc_hd__o211a_1 _16826_ (.A1(_06105_),
    .A2(_09851_),
    .B1(_09852_),
    .C1(_09812_),
    .X(_09853_));
 sky130_fd_sc_hd__a21oi_1 _16827_ (.A1(_06183_),
    .A2(_09786_),
    .B1(_09853_),
    .Y(_00534_));
 sky130_fd_sc_hd__or2_1 _16828_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .X(_09854_));
 sky130_fd_sc_hd__nand2_1 _16829_ (.A(\rbzero.wall_tracer.trackDistX[-4] ),
    .B(\rbzero.wall_tracer.stepDistX[-4] ),
    .Y(_09855_));
 sky130_fd_sc_hd__o21ai_1 _16830_ (.A1(_09847_),
    .A2(_09850_),
    .B1(_09848_),
    .Y(_09856_));
 sky130_fd_sc_hd__and3_1 _16831_ (.A(_09854_),
    .B(_09855_),
    .C(_09856_),
    .X(_09857_));
 sky130_fd_sc_hd__a21oi_1 _16832_ (.A1(_09854_),
    .A2(_09855_),
    .B1(_09856_),
    .Y(_09858_));
 sky130_fd_sc_hd__nand2_1 _16833_ (.A(_09822_),
    .B(_09347_),
    .Y(_09859_));
 sky130_fd_sc_hd__o311a_1 _16834_ (.A1(_06105_),
    .A2(_09857_),
    .A3(_09858_),
    .B1(_09812_),
    .C1(_09859_),
    .X(_09860_));
 sky130_fd_sc_hd__a21oi_1 _16835_ (.A1(_06182_),
    .A2(_09785_),
    .B1(_09860_),
    .Y(_00535_));
 sky130_fd_sc_hd__nor2_1 _16836_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_09861_));
 sky130_fd_sc_hd__nand2_1 _16837_ (.A(\rbzero.wall_tracer.trackDistX[-3] ),
    .B(\rbzero.wall_tracer.stepDistX[-3] ),
    .Y(_09862_));
 sky130_fd_sc_hd__or2b_1 _16838_ (.A(_09861_),
    .B_N(_09862_),
    .X(_09863_));
 sky130_fd_sc_hd__a21boi_1 _16839_ (.A1(_09854_),
    .A2(_09856_),
    .B1_N(_09855_),
    .Y(_09864_));
 sky130_fd_sc_hd__nor2_1 _16840_ (.A(_09863_),
    .B(_09864_),
    .Y(_09865_));
 sky130_fd_sc_hd__clkbuf_8 _16841_ (.A(_06103_),
    .X(_09866_));
 sky130_fd_sc_hd__a21o_1 _16842_ (.A1(_09863_),
    .A2(_09864_),
    .B1(_09866_),
    .X(_09867_));
 sky130_fd_sc_hd__xnor2_4 _16843_ (.A(_09355_),
    .B(_09466_),
    .Y(_09868_));
 sky130_fd_sc_hd__nand2_1 _16844_ (.A(_06104_),
    .B(_09868_),
    .Y(_09869_));
 sky130_fd_sc_hd__o21ai_1 _16845_ (.A1(_09865_),
    .A2(_09867_),
    .B1(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__mux2_1 _16846_ (.A0(\rbzero.wall_tracer.trackDistX[-3] ),
    .A1(_09870_),
    .S(_09844_),
    .X(_09871_));
 sky130_fd_sc_hd__clkbuf_1 _16847_ (.A(_09871_),
    .X(_00536_));
 sky130_fd_sc_hd__buf_4 _16848_ (.A(_06104_),
    .X(_09872_));
 sky130_fd_sc_hd__nand2_1 _16849_ (.A(_09872_),
    .B(_09593_),
    .Y(_09873_));
 sky130_fd_sc_hd__or2_1 _16850_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .X(_09874_));
 sky130_fd_sc_hd__nand2_1 _16851_ (.A(\rbzero.wall_tracer.trackDistX[-2] ),
    .B(\rbzero.wall_tracer.stepDistX[-2] ),
    .Y(_09875_));
 sky130_fd_sc_hd__o21ai_1 _16852_ (.A1(_09861_),
    .A2(_09864_),
    .B1(_09862_),
    .Y(_09876_));
 sky130_fd_sc_hd__and3_1 _16853_ (.A(_09874_),
    .B(_09875_),
    .C(_09876_),
    .X(_09877_));
 sky130_fd_sc_hd__a21oi_1 _16854_ (.A1(_09874_),
    .A2(_09875_),
    .B1(_09876_),
    .Y(_09878_));
 sky130_fd_sc_hd__buf_4 _16855_ (.A(_09782_),
    .X(_09879_));
 sky130_fd_sc_hd__o31a_1 _16856_ (.A1(_09872_),
    .A2(_09877_),
    .A3(_09878_),
    .B1(_09879_),
    .X(_09880_));
 sky130_fd_sc_hd__o2bb2a_1 _16857_ (.A1_N(_09873_),
    .A2_N(_09880_),
    .B1(\rbzero.wall_tracer.trackDistX[-2] ),
    .B2(_09879_),
    .X(_00537_));
 sky130_fd_sc_hd__nor2_1 _16858_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .Y(_09881_));
 sky130_fd_sc_hd__and2_1 _16859_ (.A(\rbzero.wall_tracer.trackDistX[-1] ),
    .B(\rbzero.wall_tracer.stepDistX[-1] ),
    .X(_09882_));
 sky130_fd_sc_hd__or2_1 _16860_ (.A(_09881_),
    .B(_09882_),
    .X(_09883_));
 sky130_fd_sc_hd__a21boi_1 _16861_ (.A1(_09874_),
    .A2(_09876_),
    .B1_N(_09875_),
    .Y(_09884_));
 sky130_fd_sc_hd__nor2_1 _16862_ (.A(_09883_),
    .B(_09884_),
    .Y(_09885_));
 sky130_fd_sc_hd__a21o_1 _16863_ (.A1(_09883_),
    .A2(_09884_),
    .B1(_09866_),
    .X(_09886_));
 sky130_fd_sc_hd__nand2_1 _16864_ (.A(_06104_),
    .B(_09721_),
    .Y(_09887_));
 sky130_fd_sc_hd__o21ai_1 _16865_ (.A1(_09885_),
    .A2(_09886_),
    .B1(_09887_),
    .Y(_09888_));
 sky130_fd_sc_hd__mux2_1 _16866_ (.A0(\rbzero.wall_tracer.trackDistX[-1] ),
    .A1(_09888_),
    .S(_09844_),
    .X(_09889_));
 sky130_fd_sc_hd__clkbuf_1 _16867_ (.A(_09889_),
    .X(_00538_));
 sky130_fd_sc_hd__clkbuf_4 _16868_ (.A(_09687_),
    .X(_09890_));
 sky130_fd_sc_hd__a31o_1 _16869_ (.A1(_08616_),
    .A2(_09607_),
    .A3(_09890_),
    .B1(_09605_),
    .X(_09891_));
 sky130_fd_sc_hd__or2b_1 _16870_ (.A(_09641_),
    .B_N(_09611_),
    .X(_09892_));
 sky130_fd_sc_hd__o2bb2a_1 _16871_ (.A1_N(_09620_),
    .A2_N(_09622_),
    .B1(_09618_),
    .B2(_09619_),
    .X(_09893_));
 sky130_fd_sc_hd__a21oi_4 _16872_ (.A1(_09639_),
    .A2(_09892_),
    .B1(_09893_),
    .Y(_09894_));
 sky130_fd_sc_hd__and3_1 _16873_ (.A(_09639_),
    .B(_09892_),
    .C(_09893_),
    .X(_09895_));
 sky130_fd_sc_hd__nor2_1 _16874_ (.A(_09894_),
    .B(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__a21o_1 _16875_ (.A1(_09623_),
    .A2(_09636_),
    .B1(_09635_),
    .X(_09897_));
 sky130_fd_sc_hd__or2b_1 _16876_ (.A(_09659_),
    .B_N(_09645_),
    .X(_09898_));
 sky130_fd_sc_hd__or2b_1 _16877_ (.A(_09660_),
    .B_N(_09643_),
    .X(_09899_));
 sky130_fd_sc_hd__nor2_1 _16878_ (.A(_08952_),
    .B(_09362_),
    .Y(_09900_));
 sky130_fd_sc_hd__xnor2_1 _16879_ (.A(_09615_),
    .B(_09900_),
    .Y(_09901_));
 sky130_fd_sc_hd__nor2_1 _16880_ (.A(_09008_),
    .B(_09490_),
    .Y(_09902_));
 sky130_fd_sc_hd__xor2_1 _16881_ (.A(_09901_),
    .B(_09902_),
    .X(_09903_));
 sky130_fd_sc_hd__nand2_1 _16882_ (.A(_09498_),
    .B(_09615_),
    .Y(_09904_));
 sky130_fd_sc_hd__o31a_1 _16883_ (.A1(_09008_),
    .A2(_09363_),
    .A3(_09616_),
    .B1(_09904_),
    .X(_09905_));
 sky130_fd_sc_hd__nor2_1 _16884_ (.A(_09903_),
    .B(_09905_),
    .Y(_09906_));
 sky130_fd_sc_hd__and2_1 _16885_ (.A(_09903_),
    .B(_09905_),
    .X(_09907_));
 sky130_fd_sc_hd__nor2_1 _16886_ (.A(_09906_),
    .B(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__or2_2 _16887_ (.A(_08159_),
    .B(_09608_),
    .X(_09909_));
 sky130_fd_sc_hd__xnor2_1 _16888_ (.A(_09908_),
    .B(_09909_),
    .Y(_09910_));
 sky130_fd_sc_hd__a21bo_1 _16889_ (.A1(_09499_),
    .A2(_09630_),
    .B1_N(_09629_),
    .X(_09911_));
 sky130_fd_sc_hd__o21ai_1 _16890_ (.A1(_09522_),
    .A2(_09649_),
    .B1(_09646_),
    .Y(_09912_));
 sky130_fd_sc_hd__o21ai_1 _16891_ (.A1(_09525_),
    .A2(_09079_),
    .B1(_09628_),
    .Y(_09913_));
 sky130_fd_sc_hd__or3_1 _16892_ (.A(_08731_),
    .B(_09079_),
    .C(_09628_),
    .X(_09914_));
 sky130_fd_sc_hd__nand2_1 _16893_ (.A(_09913_),
    .B(_09914_),
    .Y(_09915_));
 sky130_fd_sc_hd__nor2_1 _16894_ (.A(_09146_),
    .B(_09131_),
    .Y(_09916_));
 sky130_fd_sc_hd__xnor2_1 _16895_ (.A(_09915_),
    .B(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__and2_1 _16896_ (.A(_09912_),
    .B(_09917_),
    .X(_09918_));
 sky130_fd_sc_hd__or2_1 _16897_ (.A(_09912_),
    .B(_09917_),
    .X(_09919_));
 sky130_fd_sc_hd__and2b_1 _16898_ (.A_N(_09918_),
    .B(_09919_),
    .X(_09920_));
 sky130_fd_sc_hd__xnor2_1 _16899_ (.A(_09911_),
    .B(_09920_),
    .Y(_09921_));
 sky130_fd_sc_hd__nand2_1 _16900_ (.A(_09625_),
    .B(_09632_),
    .Y(_09922_));
 sky130_fd_sc_hd__a21boi_1 _16901_ (.A1(_09626_),
    .A2(_09631_),
    .B1_N(_09922_),
    .Y(_09923_));
 sky130_fd_sc_hd__xor2_1 _16902_ (.A(_09921_),
    .B(_09923_),
    .X(_09924_));
 sky130_fd_sc_hd__xnor2_1 _16903_ (.A(_09910_),
    .B(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__a21o_1 _16904_ (.A1(_09898_),
    .A2(_09899_),
    .B1(_09925_),
    .X(_09926_));
 sky130_fd_sc_hd__nand3_1 _16905_ (.A(_09898_),
    .B(_09899_),
    .C(_09925_),
    .Y(_09927_));
 sky130_fd_sc_hd__nand2_1 _16906_ (.A(_09926_),
    .B(_09927_),
    .Y(_09928_));
 sky130_fd_sc_hd__xnor2_1 _16907_ (.A(_09897_),
    .B(_09928_),
    .Y(_09929_));
 sky130_fd_sc_hd__a21o_1 _16908_ (.A1(_09650_),
    .A2(_09657_),
    .B1(_09656_),
    .X(_09930_));
 sky130_fd_sc_hd__nand2_1 _16909_ (.A(_09666_),
    .B(_09674_),
    .Y(_09931_));
 sky130_fd_sc_hd__a21bo_1 _16910_ (.A1(_09664_),
    .A2(_09675_),
    .B1_N(_09931_),
    .X(_09932_));
 sky130_fd_sc_hd__nor2_1 _16911_ (.A(_08151_),
    .B(_08580_),
    .Y(_09933_));
 sky130_fd_sc_hd__nor2_1 _16912_ (.A(_08166_),
    .B(_08382_),
    .Y(_09934_));
 sky130_fd_sc_hd__nor2_1 _16913_ (.A(_09933_),
    .B(_09934_),
    .Y(_09935_));
 sky130_fd_sc_hd__nand2_1 _16914_ (.A(_09933_),
    .B(_09934_),
    .Y(_09936_));
 sky130_fd_sc_hd__or2b_1 _16915_ (.A(_09935_),
    .B_N(_09936_),
    .X(_09937_));
 sky130_fd_sc_hd__or3_1 _16916_ (.A(_09519_),
    .B(_08620_),
    .C(_09937_),
    .X(_09938_));
 sky130_fd_sc_hd__o21ai_1 _16917_ (.A1(_09519_),
    .A2(_08620_),
    .B1(_09937_),
    .Y(_09939_));
 sky130_fd_sc_hd__and2_1 _16918_ (.A(_09938_),
    .B(_09939_),
    .X(_09940_));
 sky130_fd_sc_hd__nor2_1 _16919_ (.A(_08813_),
    .B(_09176_),
    .Y(_09941_));
 sky130_fd_sc_hd__nor2_1 _16920_ (.A(_08327_),
    .B(_09037_),
    .Y(_09942_));
 sky130_fd_sc_hd__o22a_1 _16921_ (.A1(_08327_),
    .A2(_09176_),
    .B1(_09037_),
    .B2(_08813_),
    .X(_09943_));
 sky130_fd_sc_hd__a21o_1 _16922_ (.A1(_09941_),
    .A2(_09942_),
    .B1(_09943_),
    .X(_09944_));
 sky130_fd_sc_hd__nor2_1 _16923_ (.A(_09397_),
    .B(_08497_),
    .Y(_09945_));
 sky130_fd_sc_hd__xor2_1 _16924_ (.A(_09944_),
    .B(_09945_),
    .X(_09946_));
 sky130_fd_sc_hd__or3_1 _16925_ (.A(_08373_),
    .B(_09176_),
    .C(_09651_),
    .X(_09947_));
 sky130_fd_sc_hd__a21boi_1 _16926_ (.A1(_09529_),
    .A2(_09653_),
    .B1_N(_09947_),
    .Y(_09948_));
 sky130_fd_sc_hd__nor2_1 _16927_ (.A(_09946_),
    .B(_09948_),
    .Y(_09949_));
 sky130_fd_sc_hd__nand2_1 _16928_ (.A(_09946_),
    .B(_09948_),
    .Y(_09950_));
 sky130_fd_sc_hd__and2b_1 _16929_ (.A_N(_09949_),
    .B(_09950_),
    .X(_09951_));
 sky130_fd_sc_hd__xnor2_1 _16930_ (.A(_09940_),
    .B(_09951_),
    .Y(_09952_));
 sky130_fd_sc_hd__xor2_1 _16931_ (.A(_09932_),
    .B(_09952_),
    .X(_09953_));
 sky130_fd_sc_hd__xnor2_1 _16932_ (.A(_09930_),
    .B(_09953_),
    .Y(_09954_));
 sky130_fd_sc_hd__a22o_1 _16933_ (.A1(_09557_),
    .A2(_09667_),
    .B1(_09673_),
    .B2(_09663_),
    .X(_09955_));
 sky130_fd_sc_hd__a2bb2o_1 _16934_ (.A1_N(_09679_),
    .A2_N(_09681_),
    .B1(_09682_),
    .B2(_09678_),
    .X(_09956_));
 sky130_fd_sc_hd__a21oi_1 _16935_ (.A1(_09670_),
    .A2(_09184_),
    .B1(_08516_),
    .Y(_09957_));
 sky130_fd_sc_hd__xnor2_1 _16936_ (.A(_09667_),
    .B(_09957_),
    .Y(_09958_));
 sky130_fd_sc_hd__a21o_1 _16937_ (.A1(_09044_),
    .A2(_09046_),
    .B1(_09406_),
    .X(_09959_));
 sky130_fd_sc_hd__xor2_1 _16938_ (.A(_09958_),
    .B(_09959_),
    .X(_09960_));
 sky130_fd_sc_hd__nand2_1 _16939_ (.A(_09956_),
    .B(_09960_),
    .Y(_09961_));
 sky130_fd_sc_hd__or2_1 _16940_ (.A(_09956_),
    .B(_09960_),
    .X(_09962_));
 sky130_fd_sc_hd__nand2_1 _16941_ (.A(_09961_),
    .B(_09962_),
    .Y(_09963_));
 sky130_fd_sc_hd__xnor2_2 _16942_ (.A(_09955_),
    .B(_09963_),
    .Y(_09964_));
 sky130_fd_sc_hd__nor2_1 _16943_ (.A(_09167_),
    .B(_09677_),
    .Y(_09965_));
 sky130_fd_sc_hd__nor2_1 _16944_ (.A(_08910_),
    .B(_09559_),
    .Y(_09966_));
 sky130_fd_sc_hd__xnor2_2 _16945_ (.A(_09681_),
    .B(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__xor2_2 _16946_ (.A(_09965_),
    .B(_09967_),
    .X(_09968_));
 sky130_fd_sc_hd__a2bb2oi_2 _16947_ (.A1_N(_06433_),
    .A2_N(_09691_),
    .B1(_09692_),
    .B2(_09686_),
    .Y(_09969_));
 sky130_fd_sc_hd__nand2_2 _16948_ (.A(\rbzero.wall_tracer.stepDistX[10] ),
    .B(_09045_),
    .Y(_09970_));
 sky130_fd_sc_hd__nand2_1 _16949_ (.A(\rbzero.wall_tracer.stepDistY[10] ),
    .B(_08405_),
    .Y(_09971_));
 sky130_fd_sc_hd__a21o_1 _16950_ (.A1(_09689_),
    .A2(_09971_),
    .B1(_09045_),
    .X(_09972_));
 sky130_fd_sc_hd__a21oi_1 _16951_ (.A1(_09970_),
    .A2(_09972_),
    .B1(_08950_),
    .Y(_09973_));
 sky130_fd_sc_hd__a21o_1 _16952_ (.A1(_09685_),
    .A2(_09566_),
    .B1(_09045_),
    .X(_09974_));
 sky130_fd_sc_hd__nand2_2 _16953_ (.A(\rbzero.wall_tracer.stepDistX[9] ),
    .B(_09045_),
    .Y(_09975_));
 sky130_fd_sc_hd__a21o_1 _16954_ (.A1(_09974_),
    .A2(_09975_),
    .B1(_08950_),
    .X(_09976_));
 sky130_fd_sc_hd__or3_1 _16955_ (.A(_08042_),
    .B(_08338_),
    .C(_09689_),
    .X(_09977_));
 sky130_fd_sc_hd__mux2_1 _16956_ (.A0(_08637_),
    .A1(_09977_),
    .S(_09691_),
    .X(_09978_));
 sky130_fd_sc_hd__mux2_1 _16957_ (.A0(_09973_),
    .A1(_09976_),
    .S(_09978_),
    .X(_09979_));
 sky130_fd_sc_hd__xor2_2 _16958_ (.A(_09969_),
    .B(_09979_),
    .X(_09980_));
 sky130_fd_sc_hd__xnor2_1 _16959_ (.A(_09968_),
    .B(_09980_),
    .Y(_09981_));
 sky130_fd_sc_hd__nor2_1 _16960_ (.A(_09693_),
    .B(_09695_),
    .Y(_09982_));
 sky130_fd_sc_hd__a21o_1 _16961_ (.A1(_09684_),
    .A2(_09696_),
    .B1(_09982_),
    .X(_09983_));
 sky130_fd_sc_hd__xnor2_1 _16962_ (.A(_09981_),
    .B(_09983_),
    .Y(_09984_));
 sky130_fd_sc_hd__xnor2_2 _16963_ (.A(_09964_),
    .B(_09984_),
    .Y(_09985_));
 sky130_fd_sc_hd__or2b_1 _16964_ (.A(_09697_),
    .B_N(_09699_),
    .X(_09986_));
 sky130_fd_sc_hd__a21bo_1 _16965_ (.A1(_09676_),
    .A2(_09700_),
    .B1_N(_09986_),
    .X(_09987_));
 sky130_fd_sc_hd__xnor2_1 _16966_ (.A(_09985_),
    .B(_09987_),
    .Y(_09988_));
 sky130_fd_sc_hd__xnor2_1 _16967_ (.A(_09954_),
    .B(_09988_),
    .Y(_09989_));
 sky130_fd_sc_hd__and2b_1 _16968_ (.A_N(_09701_),
    .B(_09703_),
    .X(_09990_));
 sky130_fd_sc_hd__a21oi_1 _16969_ (.A1(_09661_),
    .A2(_09704_),
    .B1(_09990_),
    .Y(_09991_));
 sky130_fd_sc_hd__or2_1 _16970_ (.A(_09989_),
    .B(_09991_),
    .X(_09992_));
 sky130_fd_sc_hd__nand2_1 _16971_ (.A(_09989_),
    .B(_09991_),
    .Y(_09993_));
 sky130_fd_sc_hd__and2_1 _16972_ (.A(_09992_),
    .B(_09993_),
    .X(_09994_));
 sky130_fd_sc_hd__xnor2_1 _16973_ (.A(_09929_),
    .B(_09994_),
    .Y(_09995_));
 sky130_fd_sc_hd__a21oi_1 _16974_ (.A1(_09642_),
    .A2(_09710_),
    .B1(_09708_),
    .Y(_09996_));
 sky130_fd_sc_hd__xor2_1 _16975_ (.A(_09995_),
    .B(_09996_),
    .X(_09997_));
 sky130_fd_sc_hd__nand2_1 _16976_ (.A(_09896_),
    .B(_09997_),
    .Y(_09998_));
 sky130_fd_sc_hd__or2_1 _16977_ (.A(_09896_),
    .B(_09997_),
    .X(_09999_));
 sky130_fd_sc_hd__nand2_1 _16978_ (.A(_09998_),
    .B(_09999_),
    .Y(_10000_));
 sky130_fd_sc_hd__o2bb2a_1 _16979_ (.A1_N(_09610_),
    .A2_N(_09713_),
    .B1(_09712_),
    .B2(_09711_),
    .X(_10001_));
 sky130_fd_sc_hd__xor2_1 _16980_ (.A(_10000_),
    .B(_10001_),
    .X(_10002_));
 sky130_fd_sc_hd__nand2_1 _16981_ (.A(_09891_),
    .B(_10002_),
    .Y(_10003_));
 sky130_fd_sc_hd__or2_1 _16982_ (.A(_09891_),
    .B(_10002_),
    .X(_10004_));
 sky130_fd_sc_hd__and2_2 _16983_ (.A(_10003_),
    .B(_10004_),
    .X(_10005_));
 sky130_fd_sc_hd__xor2_4 _16984_ (.A(_09717_),
    .B(_10005_),
    .X(_10006_));
 sky130_fd_sc_hd__inv_2 _16985_ (.A(_09720_),
    .Y(_10007_));
 sky130_fd_sc_hd__a21o_1 _16986_ (.A1(_09587_),
    .A2(_09590_),
    .B1(_09719_),
    .X(_10008_));
 sky130_fd_sc_hd__o31a_4 _16987_ (.A1(_09479_),
    .A2(_09592_),
    .A3(_10007_),
    .B1(_10008_),
    .X(_10009_));
 sky130_fd_sc_hd__xnor2_4 _16988_ (.A(_10006_),
    .B(_10009_),
    .Y(_10010_));
 sky130_fd_sc_hd__nand2_1 _16989_ (.A(_09872_),
    .B(_10010_),
    .Y(_10011_));
 sky130_fd_sc_hd__or2_1 _16990_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .X(_10012_));
 sky130_fd_sc_hd__nand2_1 _16991_ (.A(\rbzero.wall_tracer.trackDistX[0] ),
    .B(\rbzero.wall_tracer.stepDistX[0] ),
    .Y(_10013_));
 sky130_fd_sc_hd__a211oi_1 _16992_ (.A1(_10012_),
    .A2(_10013_),
    .B1(_09882_),
    .C1(_09885_),
    .Y(_10014_));
 sky130_fd_sc_hd__o211a_1 _16993_ (.A1(_09882_),
    .A2(_09885_),
    .B1(_10012_),
    .C1(_10013_),
    .X(_10015_));
 sky130_fd_sc_hd__o31a_1 _16994_ (.A1(_09872_),
    .A2(_10014_),
    .A3(_10015_),
    .B1(_09879_),
    .X(_10016_));
 sky130_fd_sc_hd__o2bb2a_1 _16995_ (.A1_N(_10011_),
    .A2_N(_10016_),
    .B1(\rbzero.wall_tracer.trackDistX[0] ),
    .B2(_09879_),
    .X(_00539_));
 sky130_fd_sc_hd__or2_1 _16996_ (.A(_10000_),
    .B(_10001_),
    .X(_10017_));
 sky130_fd_sc_hd__nand2_2 _16997_ (.A(_10017_),
    .B(_10003_),
    .Y(_10018_));
 sky130_fd_sc_hd__or2b_1 _16998_ (.A(_09928_),
    .B_N(_09897_),
    .X(_10019_));
 sky130_fd_sc_hd__o21ba_1 _16999_ (.A1(_09907_),
    .A2(_09909_),
    .B1_N(_09906_),
    .X(_10020_));
 sky130_fd_sc_hd__a21oi_1 _17000_ (.A1(_09926_),
    .A2(_10019_),
    .B1(_10020_),
    .Y(_10021_));
 sky130_fd_sc_hd__and3_1 _17001_ (.A(_09926_),
    .B(_10019_),
    .C(_10020_),
    .X(_10022_));
 sky130_fd_sc_hd__nor2_1 _17002_ (.A(_10021_),
    .B(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__nand2_1 _17003_ (.A(_09929_),
    .B(_09994_),
    .Y(_10024_));
 sky130_fd_sc_hd__nor2_1 _17004_ (.A(_09921_),
    .B(_09923_),
    .Y(_10025_));
 sky130_fd_sc_hd__a21o_1 _17005_ (.A1(_09910_),
    .A2(_09924_),
    .B1(_10025_),
    .X(_10026_));
 sky130_fd_sc_hd__or2b_1 _17006_ (.A(_09952_),
    .B_N(_09932_),
    .X(_10027_));
 sky130_fd_sc_hd__or2b_1 _17007_ (.A(_09953_),
    .B_N(_09930_),
    .X(_10028_));
 sky130_fd_sc_hd__nand2_1 _17008_ (.A(_10027_),
    .B(_10028_),
    .Y(_10029_));
 sky130_fd_sc_hd__o22a_1 _17009_ (.A1(_09146_),
    .A2(_09242_),
    .B1(_09363_),
    .B2(_09005_),
    .X(_10030_));
 sky130_fd_sc_hd__or2_1 _17010_ (.A(_09146_),
    .B(_09362_),
    .X(_10031_));
 sky130_fd_sc_hd__or3_1 _17011_ (.A(_09005_),
    .B(_09242_),
    .C(_10031_),
    .X(_10032_));
 sky130_fd_sc_hd__and2b_1 _17012_ (.A_N(_10030_),
    .B(_10032_),
    .X(_10033_));
 sky130_fd_sc_hd__nor2_1 _17013_ (.A(_08952_),
    .B(_09491_),
    .Y(_10034_));
 sky130_fd_sc_hd__xnor2_1 _17014_ (.A(_10033_),
    .B(_10034_),
    .Y(_10035_));
 sky130_fd_sc_hd__nand2_1 _17015_ (.A(_09615_),
    .B(_09900_),
    .Y(_10036_));
 sky130_fd_sc_hd__o31a_1 _17016_ (.A1(_09008_),
    .A2(_09491_),
    .A3(_09901_),
    .B1(_10036_),
    .X(_10037_));
 sky130_fd_sc_hd__xnor2_1 _17017_ (.A(_10035_),
    .B(_10037_),
    .Y(_10038_));
 sky130_fd_sc_hd__nand2_1 _17018_ (.A(_09008_),
    .B(_09890_),
    .Y(_10039_));
 sky130_fd_sc_hd__xor2_1 _17019_ (.A(_10038_),
    .B(_10039_),
    .X(_10040_));
 sky130_fd_sc_hd__o31ai_2 _17020_ (.A1(_09146_),
    .A2(_09252_),
    .A3(_09915_),
    .B1(_09914_),
    .Y(_10041_));
 sky130_fd_sc_hd__nand2_1 _17021_ (.A(_09936_),
    .B(_09938_),
    .Y(_10042_));
 sky130_fd_sc_hd__o22ai_1 _17022_ (.A1(_09519_),
    .A2(_08618_),
    .B1(_09079_),
    .B2(_09520_),
    .Y(_10043_));
 sky130_fd_sc_hd__or3_1 _17023_ (.A(_08666_),
    .B(_09079_),
    .C(_09628_),
    .X(_10044_));
 sky130_fd_sc_hd__nand2_1 _17024_ (.A(_10043_),
    .B(_10044_),
    .Y(_10045_));
 sky130_fd_sc_hd__nor2_1 _17025_ (.A(_09525_),
    .B(_09252_),
    .Y(_10046_));
 sky130_fd_sc_hd__xor2_1 _17026_ (.A(_10045_),
    .B(_10046_),
    .X(_10047_));
 sky130_fd_sc_hd__xnor2_1 _17027_ (.A(_10042_),
    .B(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__xnor2_1 _17028_ (.A(_10041_),
    .B(_10048_),
    .Y(_10049_));
 sky130_fd_sc_hd__a21oi_1 _17029_ (.A1(_09911_),
    .A2(_09919_),
    .B1(_09918_),
    .Y(_10050_));
 sky130_fd_sc_hd__nor2_1 _17030_ (.A(_10049_),
    .B(_10050_),
    .Y(_10051_));
 sky130_fd_sc_hd__and2_1 _17031_ (.A(_10049_),
    .B(_10050_),
    .X(_10052_));
 sky130_fd_sc_hd__nor2_1 _17032_ (.A(_10051_),
    .B(_10052_),
    .Y(_10053_));
 sky130_fd_sc_hd__xor2_1 _17033_ (.A(_10040_),
    .B(_10053_),
    .X(_10054_));
 sky130_fd_sc_hd__xnor2_1 _17034_ (.A(_10029_),
    .B(_10054_),
    .Y(_10055_));
 sky130_fd_sc_hd__xnor2_1 _17035_ (.A(_10026_),
    .B(_10055_),
    .Y(_10056_));
 sky130_fd_sc_hd__a21o_1 _17036_ (.A1(_09940_),
    .A2(_09950_),
    .B1(_09949_),
    .X(_10057_));
 sky130_fd_sc_hd__a21bo_1 _17037_ (.A1(_09955_),
    .A2(_09962_),
    .B1_N(_09961_),
    .X(_10058_));
 sky130_fd_sc_hd__clkbuf_4 _17038_ (.A(_08580_),
    .X(_10059_));
 sky130_fd_sc_hd__nor2_1 _17039_ (.A(_08166_),
    .B(_10059_),
    .Y(_10060_));
 sky130_fd_sc_hd__nor2_2 _17040_ (.A(_08151_),
    .B(_08399_),
    .Y(_10061_));
 sky130_fd_sc_hd__xnor2_1 _17041_ (.A(_10060_),
    .B(_10061_),
    .Y(_10062_));
 sky130_fd_sc_hd__nor2_1 _17042_ (.A(_09647_),
    .B(_08620_),
    .Y(_10063_));
 sky130_fd_sc_hd__xnor2_1 _17043_ (.A(_10062_),
    .B(_10063_),
    .Y(_10064_));
 sky130_fd_sc_hd__a21oi_1 _17044_ (.A1(_09044_),
    .A2(_09046_),
    .B1(_08813_),
    .Y(_10065_));
 sky130_fd_sc_hd__xnor2_1 _17045_ (.A(_09942_),
    .B(_10065_),
    .Y(_10066_));
 sky130_fd_sc_hd__nor2_1 _17046_ (.A(_08535_),
    .B(_09176_),
    .Y(_10067_));
 sky130_fd_sc_hd__xor2_1 _17047_ (.A(_10066_),
    .B(_10067_),
    .X(_10068_));
 sky130_fd_sc_hd__nand2_1 _17048_ (.A(_09941_),
    .B(_09942_),
    .Y(_10069_));
 sky130_fd_sc_hd__o31a_1 _17049_ (.A1(_09397_),
    .A2(_08497_),
    .A3(_09944_),
    .B1(_10069_),
    .X(_10070_));
 sky130_fd_sc_hd__nor2_1 _17050_ (.A(_10068_),
    .B(_10070_),
    .Y(_10071_));
 sky130_fd_sc_hd__nand2_1 _17051_ (.A(_10068_),
    .B(_10070_),
    .Y(_10072_));
 sky130_fd_sc_hd__and2b_1 _17052_ (.A_N(_10071_),
    .B(_10072_),
    .X(_10073_));
 sky130_fd_sc_hd__xor2_1 _17053_ (.A(_10064_),
    .B(_10073_),
    .X(_10074_));
 sky130_fd_sc_hd__xnor2_1 _17054_ (.A(_10058_),
    .B(_10074_),
    .Y(_10075_));
 sky130_fd_sc_hd__xnor2_1 _17055_ (.A(_10057_),
    .B(_10075_),
    .Y(_10076_));
 sky130_fd_sc_hd__nor2_1 _17056_ (.A(_08816_),
    .B(_09669_),
    .Y(_10077_));
 sky130_fd_sc_hd__o2bb2ai_1 _17057_ (.A1_N(_09671_),
    .A2_N(_10077_),
    .B1(_09958_),
    .B2(_09959_),
    .Y(_10078_));
 sky130_fd_sc_hd__nor2_1 _17058_ (.A(_08431_),
    .B(_09560_),
    .Y(_10079_));
 sky130_fd_sc_hd__nor2b_1 _17059_ (.A(_08910_),
    .B_N(_09680_),
    .Y(_10080_));
 sky130_fd_sc_hd__a22oi_2 _17060_ (.A1(_10079_),
    .A2(_10080_),
    .B1(_09967_),
    .B2(_09965_),
    .Y(_10081_));
 sky130_fd_sc_hd__a21oi_2 _17061_ (.A1(_09195_),
    .A2(_09421_),
    .B1(_08889_),
    .Y(_10082_));
 sky130_fd_sc_hd__xnor2_1 _17062_ (.A(_10077_),
    .B(_10082_),
    .Y(_10083_));
 sky130_fd_sc_hd__nor2_1 _17063_ (.A(_09406_),
    .B(_09186_),
    .Y(_10084_));
 sky130_fd_sc_hd__xnor2_1 _17064_ (.A(_10083_),
    .B(_10084_),
    .Y(_10085_));
 sky130_fd_sc_hd__xnor2_1 _17065_ (.A(_10081_),
    .B(_10085_),
    .Y(_10086_));
 sky130_fd_sc_hd__xor2_1 _17066_ (.A(_10078_),
    .B(_10086_),
    .X(_10087_));
 sky130_fd_sc_hd__or2_1 _17067_ (.A(_09167_),
    .B(_09560_),
    .X(_10088_));
 sky130_fd_sc_hd__a21o_1 _17068_ (.A1(_09974_),
    .A2(_09975_),
    .B1(_08431_),
    .X(_10089_));
 sky130_fd_sc_hd__xnor2_1 _17069_ (.A(_10080_),
    .B(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__xnor2_1 _17070_ (.A(_10088_),
    .B(_10090_),
    .Y(_10091_));
 sky130_fd_sc_hd__and2_1 _17071_ (.A(_09970_),
    .B(_09972_),
    .X(_10092_));
 sky130_fd_sc_hd__buf_2 _17072_ (.A(_10092_),
    .X(_10093_));
 sky130_fd_sc_hd__o211ai_1 _17073_ (.A1(_08950_),
    .A2(_10093_),
    .B1(_09977_),
    .C1(_09691_),
    .Y(_10094_));
 sky130_fd_sc_hd__o41a_1 _17074_ (.A1(_08950_),
    .A2(_08581_),
    .A3(_09691_),
    .A4(_10093_),
    .B1(_10094_),
    .X(_10095_));
 sky130_fd_sc_hd__buf_2 _17075_ (.A(_10095_),
    .X(_10096_));
 sky130_fd_sc_hd__xnor2_1 _17076_ (.A(_10091_),
    .B(_10096_),
    .Y(_10097_));
 sky130_fd_sc_hd__nor2_1 _17077_ (.A(_09969_),
    .B(_09979_),
    .Y(_10098_));
 sky130_fd_sc_hd__a21oi_1 _17078_ (.A1(_09968_),
    .A2(_09980_),
    .B1(_10098_),
    .Y(_10099_));
 sky130_fd_sc_hd__xor2_1 _17079_ (.A(_10097_),
    .B(_10099_),
    .X(_10100_));
 sky130_fd_sc_hd__xnor2_1 _17080_ (.A(_10087_),
    .B(_10100_),
    .Y(_10101_));
 sky130_fd_sc_hd__nand2_1 _17081_ (.A(_09968_),
    .B(_09980_),
    .Y(_10102_));
 sky130_fd_sc_hd__or2_1 _17082_ (.A(_09968_),
    .B(_09980_),
    .X(_10103_));
 sky130_fd_sc_hd__a32o_1 _17083_ (.A1(_10102_),
    .A2(_10103_),
    .A3(_09983_),
    .B1(_09984_),
    .B2(_09964_),
    .X(_10104_));
 sky130_fd_sc_hd__xnor2_1 _17084_ (.A(_10101_),
    .B(_10104_),
    .Y(_10105_));
 sky130_fd_sc_hd__xnor2_1 _17085_ (.A(_10076_),
    .B(_10105_),
    .Y(_10106_));
 sky130_fd_sc_hd__and2b_1 _17086_ (.A_N(_09985_),
    .B(_09987_),
    .X(_10107_));
 sky130_fd_sc_hd__a21oi_1 _17087_ (.A1(_09954_),
    .A2(_09988_),
    .B1(_10107_),
    .Y(_10108_));
 sky130_fd_sc_hd__nor2_1 _17088_ (.A(_10106_),
    .B(_10108_),
    .Y(_10109_));
 sky130_fd_sc_hd__and2_1 _17089_ (.A(_10106_),
    .B(_10108_),
    .X(_10110_));
 sky130_fd_sc_hd__nor2_1 _17090_ (.A(_10109_),
    .B(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__xnor2_1 _17091_ (.A(_10056_),
    .B(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__a21oi_1 _17092_ (.A1(_09992_),
    .A2(_10024_),
    .B1(_10112_),
    .Y(_10113_));
 sky130_fd_sc_hd__and3_1 _17093_ (.A(_09992_),
    .B(_10024_),
    .C(_10112_),
    .X(_10114_));
 sky130_fd_sc_hd__nor2_1 _17094_ (.A(_10113_),
    .B(_10114_),
    .Y(_10115_));
 sky130_fd_sc_hd__xnor2_1 _17095_ (.A(_10023_),
    .B(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__o21a_1 _17096_ (.A1(_09995_),
    .A2(_09996_),
    .B1(_09998_),
    .X(_10117_));
 sky130_fd_sc_hd__nor2_1 _17097_ (.A(_10116_),
    .B(_10117_),
    .Y(_10118_));
 sky130_fd_sc_hd__and2_1 _17098_ (.A(_10116_),
    .B(_10117_),
    .X(_10119_));
 sky130_fd_sc_hd__nor2_2 _17099_ (.A(_10118_),
    .B(_10119_),
    .Y(_10120_));
 sky130_fd_sc_hd__xnor2_4 _17100_ (.A(_09894_),
    .B(_10120_),
    .Y(_10121_));
 sky130_fd_sc_hd__xnor2_4 _17101_ (.A(_10018_),
    .B(_10121_),
    .Y(_10122_));
 sky130_fd_sc_hd__nor2_1 _17102_ (.A(_09717_),
    .B(_10005_),
    .Y(_10123_));
 sky130_fd_sc_hd__nand2_1 _17103_ (.A(_09717_),
    .B(_10005_),
    .Y(_10124_));
 sky130_fd_sc_hd__o21ai_2 _17104_ (.A1(_10123_),
    .A2(_10009_),
    .B1(_10124_),
    .Y(_10125_));
 sky130_fd_sc_hd__xor2_4 _17105_ (.A(_10122_),
    .B(_10125_),
    .X(_10126_));
 sky130_fd_sc_hd__nand2_1 _17106_ (.A(_09822_),
    .B(_10126_),
    .Y(_10127_));
 sky130_fd_sc_hd__nand2_1 _17107_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .Y(_10128_));
 sky130_fd_sc_hd__or2_1 _17108_ (.A(\rbzero.wall_tracer.trackDistX[1] ),
    .B(\rbzero.wall_tracer.stepDistX[1] ),
    .X(_10129_));
 sky130_fd_sc_hd__a21o_1 _17109_ (.A1(\rbzero.wall_tracer.trackDistX[0] ),
    .A2(\rbzero.wall_tracer.stepDistX[0] ),
    .B1(_10015_),
    .X(_10130_));
 sky130_fd_sc_hd__and3_1 _17110_ (.A(_10128_),
    .B(_10129_),
    .C(_10130_),
    .X(_10131_));
 sky130_fd_sc_hd__a21o_1 _17111_ (.A1(_10128_),
    .A2(_10129_),
    .B1(_10130_),
    .X(_10132_));
 sky130_fd_sc_hd__or3b_1 _17112_ (.A(_09866_),
    .B(_10131_),
    .C_N(_10132_),
    .X(_10133_));
 sky130_fd_sc_hd__and3_1 _17113_ (.A(_09782_),
    .B(_10127_),
    .C(_10133_),
    .X(_10134_));
 sky130_fd_sc_hd__a21oi_1 _17114_ (.A1(_06202_),
    .A2(_09785_),
    .B1(_10134_),
    .Y(_00540_));
 sky130_fd_sc_hd__nand2_1 _17115_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .Y(_10135_));
 sky130_fd_sc_hd__or2_1 _17116_ (.A(\rbzero.wall_tracer.trackDistX[2] ),
    .B(\rbzero.wall_tracer.stepDistX[2] ),
    .X(_10136_));
 sky130_fd_sc_hd__inv_2 _17117_ (.A(_10128_),
    .Y(_10137_));
 sky130_fd_sc_hd__a211o_1 _17118_ (.A1(_10135_),
    .A2(_10136_),
    .B1(_10137_),
    .C1(_10131_),
    .X(_10138_));
 sky130_fd_sc_hd__o211ai_2 _17119_ (.A1(_10137_),
    .A2(_10131_),
    .B1(_10135_),
    .C1(_10136_),
    .Y(_10139_));
 sky130_fd_sc_hd__nand2_1 _17120_ (.A(_10138_),
    .B(_10139_),
    .Y(_10140_));
 sky130_fd_sc_hd__nand2_1 _17121_ (.A(_10029_),
    .B(_10054_),
    .Y(_10141_));
 sky130_fd_sc_hd__or2b_1 _17122_ (.A(_10055_),
    .B_N(_10026_),
    .X(_10142_));
 sky130_fd_sc_hd__o22a_1 _17123_ (.A1(_10035_),
    .A2(_10037_),
    .B1(_10038_),
    .B2(_10039_),
    .X(_10143_));
 sky130_fd_sc_hd__a21oi_1 _17124_ (.A1(_10141_),
    .A2(_10142_),
    .B1(_10143_),
    .Y(_10144_));
 sky130_fd_sc_hd__and3_1 _17125_ (.A(_10141_),
    .B(_10142_),
    .C(_10143_),
    .X(_10145_));
 sky130_fd_sc_hd__nor2_1 _17126_ (.A(_10144_),
    .B(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__a21o_1 _17127_ (.A1(_10040_),
    .A2(_10053_),
    .B1(_10051_),
    .X(_10147_));
 sky130_fd_sc_hd__or2b_1 _17128_ (.A(_10075_),
    .B_N(_10057_),
    .X(_10148_));
 sky130_fd_sc_hd__a21bo_1 _17129_ (.A1(_10058_),
    .A2(_10074_),
    .B1_N(_10148_),
    .X(_10149_));
 sky130_fd_sc_hd__nor2_1 _17130_ (.A(_09525_),
    .B(_09242_),
    .Y(_10150_));
 sky130_fd_sc_hd__xnor2_1 _17131_ (.A(_10031_),
    .B(_10150_),
    .Y(_10151_));
 sky130_fd_sc_hd__nor2_1 _17132_ (.A(_09005_),
    .B(_09491_),
    .Y(_10152_));
 sky130_fd_sc_hd__nand2_1 _17133_ (.A(_10151_),
    .B(_10152_),
    .Y(_10153_));
 sky130_fd_sc_hd__or2_1 _17134_ (.A(_10151_),
    .B(_10152_),
    .X(_10154_));
 sky130_fd_sc_hd__nand2_1 _17135_ (.A(_10153_),
    .B(_10154_),
    .Y(_10155_));
 sky130_fd_sc_hd__o31a_1 _17136_ (.A1(_08952_),
    .A2(_09491_),
    .A3(_10030_),
    .B1(_10032_),
    .X(_10156_));
 sky130_fd_sc_hd__xor2_1 _17137_ (.A(_10155_),
    .B(_10156_),
    .X(_10157_));
 sky130_fd_sc_hd__and2_1 _17138_ (.A(_08952_),
    .B(_09890_),
    .X(_10158_));
 sky130_fd_sc_hd__xor2_1 _17139_ (.A(_10157_),
    .B(_10158_),
    .X(_10159_));
 sky130_fd_sc_hd__a21bo_1 _17140_ (.A1(_10043_),
    .A2(_10046_),
    .B1_N(_10044_),
    .X(_10160_));
 sky130_fd_sc_hd__o22ai_1 _17141_ (.A1(_08382_),
    .A2(_08618_),
    .B1(_09079_),
    .B2(_08666_),
    .Y(_10161_));
 sky130_fd_sc_hd__or4_1 _17142_ (.A(_08666_),
    .B(_08382_),
    .C(_08617_),
    .D(_09079_),
    .X(_10162_));
 sky130_fd_sc_hd__nand2_1 _17143_ (.A(_10161_),
    .B(_10162_),
    .Y(_10163_));
 sky130_fd_sc_hd__nor2_1 _17144_ (.A(_09520_),
    .B(_09252_),
    .Y(_10164_));
 sky130_fd_sc_hd__xor2_1 _17145_ (.A(_10163_),
    .B(_10164_),
    .X(_10165_));
 sky130_fd_sc_hd__nand2_1 _17146_ (.A(_10060_),
    .B(_10061_),
    .Y(_10166_));
 sky130_fd_sc_hd__o31ai_1 _17147_ (.A1(_09647_),
    .A2(_08620_),
    .A3(_10062_),
    .B1(_10166_),
    .Y(_10167_));
 sky130_fd_sc_hd__and2b_1 _17148_ (.A_N(_10165_),
    .B(_10167_),
    .X(_10168_));
 sky130_fd_sc_hd__and2b_1 _17149_ (.A_N(_10167_),
    .B(_10165_),
    .X(_10169_));
 sky130_fd_sc_hd__nor2_1 _17150_ (.A(_10168_),
    .B(_10169_),
    .Y(_10170_));
 sky130_fd_sc_hd__xnor2_1 _17151_ (.A(_10160_),
    .B(_10170_),
    .Y(_10171_));
 sky130_fd_sc_hd__a21oi_1 _17152_ (.A1(_09936_),
    .A2(_09938_),
    .B1(_10047_),
    .Y(_10172_));
 sky130_fd_sc_hd__a21oi_1 _17153_ (.A1(_10041_),
    .A2(_10048_),
    .B1(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__nor2_1 _17154_ (.A(_10171_),
    .B(_10173_),
    .Y(_10174_));
 sky130_fd_sc_hd__and2_1 _17155_ (.A(_10171_),
    .B(_10173_),
    .X(_10175_));
 sky130_fd_sc_hd__nor2_1 _17156_ (.A(_10174_),
    .B(_10175_),
    .Y(_10176_));
 sky130_fd_sc_hd__xor2_1 _17157_ (.A(_10159_),
    .B(_10176_),
    .X(_10177_));
 sky130_fd_sc_hd__xnor2_1 _17158_ (.A(_10149_),
    .B(_10177_),
    .Y(_10178_));
 sky130_fd_sc_hd__xnor2_1 _17159_ (.A(_10147_),
    .B(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__a21o_1 _17160_ (.A1(_10064_),
    .A2(_10072_),
    .B1(_10071_),
    .X(_10180_));
 sky130_fd_sc_hd__and2b_1 _17161_ (.A_N(_10081_),
    .B(_10085_),
    .X(_10181_));
 sky130_fd_sc_hd__a21oi_1 _17162_ (.A1(_10078_),
    .A2(_10086_),
    .B1(_10181_),
    .Y(_10182_));
 sky130_fd_sc_hd__nor2_1 _17163_ (.A(_08338_),
    .B(_08499_),
    .Y(_10183_));
 sky130_fd_sc_hd__o22a_1 _17164_ (.A1(_08165_),
    .A2(_08399_),
    .B1(_08499_),
    .B2(_08151_),
    .X(_10184_));
 sky130_fd_sc_hd__a41o_1 _17165_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_08421_),
    .A3(_10183_),
    .A4(_10061_),
    .B1(_10184_),
    .X(_10185_));
 sky130_fd_sc_hd__or3_1 _17166_ (.A(_10059_),
    .B(_08553_),
    .C(_10185_),
    .X(_10186_));
 sky130_fd_sc_hd__o21ai_1 _17167_ (.A1(_10059_),
    .A2(_08620_),
    .B1(_10185_),
    .Y(_10187_));
 sky130_fd_sc_hd__and2_1 _17168_ (.A(_10186_),
    .B(_10187_),
    .X(_10188_));
 sky130_fd_sc_hd__a21oi_1 _17169_ (.A1(_09044_),
    .A2(_09046_),
    .B1(_09528_),
    .Y(_10189_));
 sky130_fd_sc_hd__a21oi_2 _17170_ (.A1(_09670_),
    .A2(_09184_),
    .B1(_08813_),
    .Y(_10190_));
 sky130_fd_sc_hd__xnor2_1 _17171_ (.A(_10189_),
    .B(_10190_),
    .Y(_10191_));
 sky130_fd_sc_hd__or2_1 _17172_ (.A(_08535_),
    .B(_09037_),
    .X(_10192_));
 sky130_fd_sc_hd__xnor2_1 _17173_ (.A(_10191_),
    .B(_10192_),
    .Y(_10193_));
 sky130_fd_sc_hd__nand2_1 _17174_ (.A(_09942_),
    .B(_10065_),
    .Y(_10194_));
 sky130_fd_sc_hd__o31a_1 _17175_ (.A1(_09397_),
    .A2(_09176_),
    .A3(_10066_),
    .B1(_10194_),
    .X(_10195_));
 sky130_fd_sc_hd__nor2_1 _17176_ (.A(_10193_),
    .B(_10195_),
    .Y(_10196_));
 sky130_fd_sc_hd__nand2_1 _17177_ (.A(_10193_),
    .B(_10195_),
    .Y(_10197_));
 sky130_fd_sc_hd__and2b_1 _17178_ (.A_N(_10196_),
    .B(_10197_),
    .X(_10198_));
 sky130_fd_sc_hd__xor2_1 _17179_ (.A(_10188_),
    .B(_10198_),
    .X(_10199_));
 sky130_fd_sc_hd__xnor2_1 _17180_ (.A(_10182_),
    .B(_10199_),
    .Y(_10200_));
 sky130_fd_sc_hd__xor2_1 _17181_ (.A(_10180_),
    .B(_10200_),
    .X(_10201_));
 sky130_fd_sc_hd__nand2_1 _17182_ (.A(_10077_),
    .B(_10082_),
    .Y(_10202_));
 sky130_fd_sc_hd__o31ai_2 _17183_ (.A1(_09542_),
    .A2(_09186_),
    .A3(_10083_),
    .B1(_10202_),
    .Y(_10203_));
 sky130_fd_sc_hd__a21o_1 _17184_ (.A1(_09974_),
    .A2(_09975_),
    .B1(_08910_),
    .X(_10204_));
 sky130_fd_sc_hd__and2b_1 _17185_ (.A_N(_10080_),
    .B(_10089_),
    .X(_10205_));
 sky130_fd_sc_hd__o22a_1 _17186_ (.A1(_09681_),
    .A2(_10204_),
    .B1(_10205_),
    .B2(_10088_),
    .X(_10206_));
 sky130_fd_sc_hd__or3b_1 _17187_ (.A(_08816_),
    .B(_09560_),
    .C_N(_10082_),
    .X(_10207_));
 sky130_fd_sc_hd__o22ai_1 _17188_ (.A1(_08816_),
    .A2(_09677_),
    .B1(_09560_),
    .B2(_08889_),
    .Y(_10208_));
 sky130_fd_sc_hd__nand2_1 _17189_ (.A(_10207_),
    .B(_10208_),
    .Y(_10209_));
 sky130_fd_sc_hd__nor2_1 _17190_ (.A(_09406_),
    .B(_09669_),
    .Y(_10210_));
 sky130_fd_sc_hd__xnor2_1 _17191_ (.A(_10209_),
    .B(_10210_),
    .Y(_10211_));
 sky130_fd_sc_hd__xnor2_1 _17192_ (.A(_10206_),
    .B(_10211_),
    .Y(_10212_));
 sky130_fd_sc_hd__xor2_1 _17193_ (.A(_10203_),
    .B(_10212_),
    .X(_10213_));
 sky130_fd_sc_hd__nand2_1 _17194_ (.A(_06263_),
    .B(_09426_),
    .Y(_10214_));
 sky130_fd_sc_hd__a21boi_4 _17195_ (.A1(\rbzero.wall_tracer.stepDistX[8] ),
    .A2(_09045_),
    .B1_N(_10214_),
    .Y(_10215_));
 sky130_fd_sc_hd__nor2_1 _17196_ (.A(_09167_),
    .B(_10215_),
    .Y(_10216_));
 sky130_fd_sc_hd__a21oi_1 _17197_ (.A1(_09970_),
    .A2(_09972_),
    .B1(_08431_),
    .Y(_10217_));
 sky130_fd_sc_hd__xnor2_1 _17198_ (.A(_10204_),
    .B(_10217_),
    .Y(_10218_));
 sky130_fd_sc_hd__xor2_2 _17199_ (.A(_10216_),
    .B(_10218_),
    .X(_10219_));
 sky130_fd_sc_hd__xor2_1 _17200_ (.A(_10096_),
    .B(_10219_),
    .X(_10220_));
 sky130_fd_sc_hd__nor3b_4 _17201_ (.A(_08581_),
    .B(_09691_),
    .C_N(_09973_),
    .Y(_10221_));
 sky130_fd_sc_hd__a21o_1 _17202_ (.A1(_10091_),
    .A2(_10096_),
    .B1(_10221_),
    .X(_10222_));
 sky130_fd_sc_hd__xor2_1 _17203_ (.A(_10220_),
    .B(_10222_),
    .X(_10223_));
 sky130_fd_sc_hd__xnor2_1 _17204_ (.A(_10213_),
    .B(_10223_),
    .Y(_10224_));
 sky130_fd_sc_hd__nor2_1 _17205_ (.A(_10097_),
    .B(_10099_),
    .Y(_10225_));
 sky130_fd_sc_hd__a21o_1 _17206_ (.A1(_10087_),
    .A2(_10100_),
    .B1(_10225_),
    .X(_10226_));
 sky130_fd_sc_hd__xnor2_1 _17207_ (.A(_10224_),
    .B(_10226_),
    .Y(_10227_));
 sky130_fd_sc_hd__xnor2_1 _17208_ (.A(_10201_),
    .B(_10227_),
    .Y(_10228_));
 sky130_fd_sc_hd__and2b_1 _17209_ (.A_N(_10101_),
    .B(_10104_),
    .X(_10229_));
 sky130_fd_sc_hd__a21oi_1 _17210_ (.A1(_10076_),
    .A2(_10105_),
    .B1(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__nor2_1 _17211_ (.A(_10228_),
    .B(_10230_),
    .Y(_10231_));
 sky130_fd_sc_hd__and2_1 _17212_ (.A(_10228_),
    .B(_10230_),
    .X(_10232_));
 sky130_fd_sc_hd__nor2_1 _17213_ (.A(_10231_),
    .B(_10232_),
    .Y(_10233_));
 sky130_fd_sc_hd__xnor2_1 _17214_ (.A(_10179_),
    .B(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__a21oi_1 _17215_ (.A1(_10056_),
    .A2(_10111_),
    .B1(_10109_),
    .Y(_10235_));
 sky130_fd_sc_hd__nor2_1 _17216_ (.A(_10234_),
    .B(_10235_),
    .Y(_10236_));
 sky130_fd_sc_hd__and2_1 _17217_ (.A(_10234_),
    .B(_10235_),
    .X(_10237_));
 sky130_fd_sc_hd__nor2_1 _17218_ (.A(_10236_),
    .B(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__xnor2_1 _17219_ (.A(_10146_),
    .B(_10238_),
    .Y(_10239_));
 sky130_fd_sc_hd__a21oi_1 _17220_ (.A1(_10023_),
    .A2(_10115_),
    .B1(_10113_),
    .Y(_10240_));
 sky130_fd_sc_hd__xor2_1 _17221_ (.A(_10239_),
    .B(_10240_),
    .X(_10241_));
 sky130_fd_sc_hd__nand2_1 _17222_ (.A(_10021_),
    .B(_10241_),
    .Y(_10242_));
 sky130_fd_sc_hd__or2_1 _17223_ (.A(_10021_),
    .B(_10241_),
    .X(_10243_));
 sky130_fd_sc_hd__nand2_1 _17224_ (.A(_10242_),
    .B(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__a21oi_1 _17225_ (.A1(_09894_),
    .A2(_10120_),
    .B1(_10118_),
    .Y(_10245_));
 sky130_fd_sc_hd__or2_1 _17226_ (.A(_10244_),
    .B(_10245_),
    .X(_10246_));
 sky130_fd_sc_hd__nand2_1 _17227_ (.A(_10244_),
    .B(_10245_),
    .Y(_10247_));
 sky130_fd_sc_hd__and2_1 _17228_ (.A(_10246_),
    .B(_10247_),
    .X(_10248_));
 sky130_fd_sc_hd__nand2_1 _17229_ (.A(_10006_),
    .B(_10122_),
    .Y(_10249_));
 sky130_fd_sc_hd__a21o_1 _17230_ (.A1(_10017_),
    .A2(_10003_),
    .B1(_10121_),
    .X(_10250_));
 sky130_fd_sc_hd__and3_1 _17231_ (.A(_10017_),
    .B(_10003_),
    .C(_10121_),
    .X(_10251_));
 sky130_fd_sc_hd__a21o_1 _17232_ (.A1(_10124_),
    .A2(_10250_),
    .B1(_10251_),
    .X(_10252_));
 sky130_fd_sc_hd__o21ai_2 _17233_ (.A1(_10009_),
    .A2(_10249_),
    .B1(_10252_),
    .Y(_10253_));
 sky130_fd_sc_hd__nand2_1 _17234_ (.A(_10248_),
    .B(_10253_),
    .Y(_10254_));
 sky130_fd_sc_hd__inv_2 _17235_ (.A(_10248_),
    .Y(_10255_));
 sky130_fd_sc_hd__o21a_1 _17236_ (.A1(_10009_),
    .A2(_10249_),
    .B1(_10252_),
    .X(_10256_));
 sky130_fd_sc_hd__nand2_1 _17237_ (.A(_10255_),
    .B(_10256_),
    .Y(_10257_));
 sky130_fd_sc_hd__and2_2 _17238_ (.A(_10254_),
    .B(_10257_),
    .X(_10258_));
 sky130_fd_sc_hd__nand2_1 _17239_ (.A(_09822_),
    .B(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__o211a_1 _17240_ (.A1(_06105_),
    .A2(_10140_),
    .B1(_10259_),
    .C1(_09812_),
    .X(_10260_));
 sky130_fd_sc_hd__a21oi_1 _17241_ (.A1(_06172_),
    .A2(_09785_),
    .B1(_10260_),
    .Y(_00541_));
 sky130_fd_sc_hd__and2_1 _17242_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .X(_10261_));
 sky130_fd_sc_hd__nor2_1 _17243_ (.A(\rbzero.wall_tracer.trackDistX[3] ),
    .B(\rbzero.wall_tracer.stepDistX[3] ),
    .Y(_10262_));
 sky130_fd_sc_hd__o211a_1 _17244_ (.A1(_10261_),
    .A2(_10262_),
    .B1(_10135_),
    .C1(_10139_),
    .X(_10263_));
 sky130_fd_sc_hd__a211oi_2 _17245_ (.A1(_10135_),
    .A2(_10139_),
    .B1(_10261_),
    .C1(_10262_),
    .Y(_10264_));
 sky130_fd_sc_hd__or2_1 _17246_ (.A(_10239_),
    .B(_10240_),
    .X(_10265_));
 sky130_fd_sc_hd__nand2_1 _17247_ (.A(_10149_),
    .B(_10177_),
    .Y(_10266_));
 sky130_fd_sc_hd__or2b_1 _17248_ (.A(_10178_),
    .B_N(_10147_),
    .X(_10267_));
 sky130_fd_sc_hd__o2bb2a_1 _17249_ (.A1_N(_10157_),
    .A2_N(_10158_),
    .B1(_10155_),
    .B2(_10156_),
    .X(_10268_));
 sky130_fd_sc_hd__a21oi_1 _17250_ (.A1(_10266_),
    .A2(_10267_),
    .B1(_10268_),
    .Y(_10269_));
 sky130_fd_sc_hd__and3_1 _17251_ (.A(_10266_),
    .B(_10267_),
    .C(_10268_),
    .X(_10270_));
 sky130_fd_sc_hd__nor2_1 _17252_ (.A(_10269_),
    .B(_10270_),
    .Y(_10271_));
 sky130_fd_sc_hd__a21o_1 _17253_ (.A1(_10159_),
    .A2(_10176_),
    .B1(_10174_),
    .X(_10272_));
 sky130_fd_sc_hd__or2b_1 _17254_ (.A(_10182_),
    .B_N(_10199_),
    .X(_10273_));
 sky130_fd_sc_hd__a21bo_1 _17255_ (.A1(_10180_),
    .A2(_10200_),
    .B1_N(_10273_),
    .X(_10274_));
 sky130_fd_sc_hd__nor2_1 _17256_ (.A(_09520_),
    .B(_09362_),
    .Y(_10275_));
 sky130_fd_sc_hd__or2_1 _17257_ (.A(_09520_),
    .B(_09242_),
    .X(_10276_));
 sky130_fd_sc_hd__o21a_1 _17258_ (.A1(_09525_),
    .A2(_09362_),
    .B1(_10276_),
    .X(_10277_));
 sky130_fd_sc_hd__a21oi_1 _17259_ (.A1(_10150_),
    .A2(_10275_),
    .B1(_10277_),
    .Y(_10278_));
 sky130_fd_sc_hd__nor2_1 _17260_ (.A(_09146_),
    .B(_09490_),
    .Y(_10279_));
 sky130_fd_sc_hd__and2_1 _17261_ (.A(_10278_),
    .B(_10279_),
    .X(_10280_));
 sky130_fd_sc_hd__nor2_1 _17262_ (.A(_10278_),
    .B(_10279_),
    .Y(_10281_));
 sky130_fd_sc_hd__or2_1 _17263_ (.A(_10280_),
    .B(_10281_),
    .X(_10282_));
 sky130_fd_sc_hd__o31a_1 _17264_ (.A1(_09525_),
    .A2(_09243_),
    .A3(_10031_),
    .B1(_10153_),
    .X(_10283_));
 sky130_fd_sc_hd__xor2_1 _17265_ (.A(_10282_),
    .B(_10283_),
    .X(_10284_));
 sky130_fd_sc_hd__and2_1 _17266_ (.A(_09005_),
    .B(_09687_),
    .X(_10285_));
 sky130_fd_sc_hd__xor2_1 _17267_ (.A(_10284_),
    .B(_10285_),
    .X(_10286_));
 sky130_fd_sc_hd__a21bo_1 _17268_ (.A1(_10161_),
    .A2(_10164_),
    .B1_N(_10162_),
    .X(_10287_));
 sky130_fd_sc_hd__nand2_2 _17269_ (.A(\rbzero.wall_tracer.visualWallDist[2] ),
    .B(_08421_),
    .Y(_10288_));
 sky130_fd_sc_hd__or2_1 _17270_ (.A(_10288_),
    .B(_08428_),
    .X(_10289_));
 sky130_fd_sc_hd__or3_1 _17271_ (.A(_08152_),
    .B(_08399_),
    .C(_10289_),
    .X(_10290_));
 sky130_fd_sc_hd__o22ai_1 _17272_ (.A1(_08580_),
    .A2(_08618_),
    .B1(_09079_),
    .B2(_08382_),
    .Y(_10291_));
 sky130_fd_sc_hd__or4_1 _17273_ (.A(_08580_),
    .B(_08382_),
    .C(_08617_),
    .D(_09076_),
    .X(_10292_));
 sky130_fd_sc_hd__nand2_1 _17274_ (.A(_10291_),
    .B(_10292_),
    .Y(_10293_));
 sky130_fd_sc_hd__nor2_1 _17275_ (.A(_08666_),
    .B(_09131_),
    .Y(_10294_));
 sky130_fd_sc_hd__xor2_1 _17276_ (.A(_10293_),
    .B(_10294_),
    .X(_10295_));
 sky130_fd_sc_hd__a21oi_1 _17277_ (.A1(_10290_),
    .A2(_10186_),
    .B1(_10295_),
    .Y(_10296_));
 sky130_fd_sc_hd__and3_1 _17278_ (.A(_10290_),
    .B(_10186_),
    .C(_10295_),
    .X(_10297_));
 sky130_fd_sc_hd__nor2_1 _17279_ (.A(_10296_),
    .B(_10297_),
    .Y(_10298_));
 sky130_fd_sc_hd__xnor2_1 _17280_ (.A(_10287_),
    .B(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__a21oi_1 _17281_ (.A1(_10160_),
    .A2(_10170_),
    .B1(_10168_),
    .Y(_10300_));
 sky130_fd_sc_hd__nor2_1 _17282_ (.A(_10299_),
    .B(_10300_),
    .Y(_10301_));
 sky130_fd_sc_hd__and2_1 _17283_ (.A(_10299_),
    .B(_10300_),
    .X(_10302_));
 sky130_fd_sc_hd__nor2_1 _17284_ (.A(_10301_),
    .B(_10302_),
    .Y(_10303_));
 sky130_fd_sc_hd__xor2_1 _17285_ (.A(_10286_),
    .B(_10303_),
    .X(_10304_));
 sky130_fd_sc_hd__nand2_1 _17286_ (.A(_10274_),
    .B(_10304_),
    .Y(_10305_));
 sky130_fd_sc_hd__or2_1 _17287_ (.A(_10274_),
    .B(_10304_),
    .X(_10306_));
 sky130_fd_sc_hd__nand2_1 _17288_ (.A(_10305_),
    .B(_10306_),
    .Y(_10307_));
 sky130_fd_sc_hd__xnor2_1 _17289_ (.A(_10272_),
    .B(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__a21o_1 _17290_ (.A1(_10188_),
    .A2(_10197_),
    .B1(_10196_),
    .X(_10309_));
 sky130_fd_sc_hd__and2b_1 _17291_ (.A_N(_10206_),
    .B(_10211_),
    .X(_10310_));
 sky130_fd_sc_hd__a21oi_1 _17292_ (.A1(_10203_),
    .A2(_10212_),
    .B1(_10310_),
    .Y(_10311_));
 sky130_fd_sc_hd__and3_1 _17293_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08475_),
    .C(_08445_),
    .X(_10312_));
 sky130_fd_sc_hd__xor2_1 _17294_ (.A(_10289_),
    .B(_10312_),
    .X(_10313_));
 sky130_fd_sc_hd__or3_1 _17295_ (.A(_08399_),
    .B(_08553_),
    .C(_10313_),
    .X(_10314_));
 sky130_fd_sc_hd__buf_2 _17296_ (.A(_08399_),
    .X(_10315_));
 sky130_fd_sc_hd__o21ai_1 _17297_ (.A1(_10315_),
    .A2(_08620_),
    .B1(_10313_),
    .Y(_10316_));
 sky130_fd_sc_hd__and2_1 _17298_ (.A(_10314_),
    .B(_10316_),
    .X(_10317_));
 sky130_fd_sc_hd__nor2_1 _17299_ (.A(_09528_),
    .B(_09669_),
    .Y(_10318_));
 sky130_fd_sc_hd__o22a_1 _17300_ (.A1(_09528_),
    .A2(_09186_),
    .B1(_09669_),
    .B2(_08814_),
    .X(_10319_));
 sky130_fd_sc_hd__a21oi_1 _17301_ (.A1(_10190_),
    .A2(_10318_),
    .B1(_10319_),
    .Y(_10320_));
 sky130_fd_sc_hd__a21oi_2 _17302_ (.A1(_09662_),
    .A2(_09046_),
    .B1(_09397_),
    .Y(_10321_));
 sky130_fd_sc_hd__xnor2_1 _17303_ (.A(_10320_),
    .B(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__nand2_1 _17304_ (.A(_10189_),
    .B(_10190_),
    .Y(_10323_));
 sky130_fd_sc_hd__o31a_1 _17305_ (.A1(_09397_),
    .A2(_09037_),
    .A3(_10191_),
    .B1(_10323_),
    .X(_10324_));
 sky130_fd_sc_hd__xor2_1 _17306_ (.A(_10322_),
    .B(_10324_),
    .X(_10325_));
 sky130_fd_sc_hd__xnor2_1 _17307_ (.A(_10317_),
    .B(_10325_),
    .Y(_10326_));
 sky130_fd_sc_hd__xnor2_1 _17308_ (.A(_10311_),
    .B(_10326_),
    .Y(_10327_));
 sky130_fd_sc_hd__xnor2_1 _17309_ (.A(_10309_),
    .B(_10327_),
    .Y(_10328_));
 sky130_fd_sc_hd__a21bo_1 _17310_ (.A1(_10208_),
    .A2(_10210_),
    .B1_N(_10207_),
    .X(_10329_));
 sky130_fd_sc_hd__and2_1 _17311_ (.A(_09974_),
    .B(_09975_),
    .X(_10330_));
 sky130_fd_sc_hd__a211o_1 _17312_ (.A1(_09970_),
    .A2(_09972_),
    .B1(_08410_),
    .C1(_08390_),
    .X(_10331_));
 sky130_fd_sc_hd__a2bb2o_1 _17313_ (.A1_N(_10330_),
    .A2_N(_10331_),
    .B1(_10218_),
    .B2(_10216_),
    .X(_10332_));
 sky130_fd_sc_hd__nor2_1 _17314_ (.A(_08816_),
    .B(_09559_),
    .Y(_10333_));
 sky130_fd_sc_hd__and2b_1 _17315_ (.A_N(_08889_),
    .B(_09680_),
    .X(_10334_));
 sky130_fd_sc_hd__xnor2_1 _17316_ (.A(_10333_),
    .B(_10334_),
    .Y(_10335_));
 sky130_fd_sc_hd__nor2_1 _17317_ (.A(_09406_),
    .B(_09677_),
    .Y(_10336_));
 sky130_fd_sc_hd__xnor2_1 _17318_ (.A(_10335_),
    .B(_10336_),
    .Y(_10337_));
 sky130_fd_sc_hd__xnor2_1 _17319_ (.A(_10332_),
    .B(_10337_),
    .Y(_10338_));
 sky130_fd_sc_hd__xnor2_1 _17320_ (.A(_10329_),
    .B(_10338_),
    .Y(_10339_));
 sky130_fd_sc_hd__and2_1 _17321_ (.A(_08410_),
    .B(_08390_),
    .X(_10340_));
 sky130_fd_sc_hd__or3b_1 _17322_ (.A(_10340_),
    .B(_10092_),
    .C_N(_10331_),
    .X(_10341_));
 sky130_fd_sc_hd__clkbuf_2 _17323_ (.A(_10341_),
    .X(_10342_));
 sky130_fd_sc_hd__nor2_1 _17324_ (.A(_09167_),
    .B(_10330_),
    .Y(_10343_));
 sky130_fd_sc_hd__xnor2_1 _17325_ (.A(_10342_),
    .B(_10343_),
    .Y(_10344_));
 sky130_fd_sc_hd__xnor2_1 _17326_ (.A(_10096_),
    .B(_10344_),
    .Y(_10345_));
 sky130_fd_sc_hd__a21oi_1 _17327_ (.A1(_10096_),
    .A2(_10219_),
    .B1(_10221_),
    .Y(_10346_));
 sky130_fd_sc_hd__xor2_1 _17328_ (.A(_10345_),
    .B(_10346_),
    .X(_10347_));
 sky130_fd_sc_hd__xnor2_1 _17329_ (.A(_10339_),
    .B(_10347_),
    .Y(_10348_));
 sky130_fd_sc_hd__nand2_1 _17330_ (.A(_10220_),
    .B(_10222_),
    .Y(_10349_));
 sky130_fd_sc_hd__a21bo_1 _17331_ (.A1(_10213_),
    .A2(_10223_),
    .B1_N(_10349_),
    .X(_10350_));
 sky130_fd_sc_hd__xnor2_1 _17332_ (.A(_10348_),
    .B(_10350_),
    .Y(_10351_));
 sky130_fd_sc_hd__xnor2_1 _17333_ (.A(_10328_),
    .B(_10351_),
    .Y(_10352_));
 sky130_fd_sc_hd__and2b_1 _17334_ (.A_N(_10224_),
    .B(_10226_),
    .X(_10353_));
 sky130_fd_sc_hd__a21oi_1 _17335_ (.A1(_10201_),
    .A2(_10227_),
    .B1(_10353_),
    .Y(_10354_));
 sky130_fd_sc_hd__nor2_1 _17336_ (.A(_10352_),
    .B(_10354_),
    .Y(_10355_));
 sky130_fd_sc_hd__and2_1 _17337_ (.A(_10352_),
    .B(_10354_),
    .X(_10356_));
 sky130_fd_sc_hd__nor2_1 _17338_ (.A(_10355_),
    .B(_10356_),
    .Y(_10357_));
 sky130_fd_sc_hd__xnor2_1 _17339_ (.A(_10308_),
    .B(_10357_),
    .Y(_10358_));
 sky130_fd_sc_hd__a21oi_1 _17340_ (.A1(_10179_),
    .A2(_10233_),
    .B1(_10231_),
    .Y(_10359_));
 sky130_fd_sc_hd__xor2_1 _17341_ (.A(_10358_),
    .B(_10359_),
    .X(_10360_));
 sky130_fd_sc_hd__nand2_1 _17342_ (.A(_10271_),
    .B(_10360_),
    .Y(_10361_));
 sky130_fd_sc_hd__or2_1 _17343_ (.A(_10271_),
    .B(_10360_),
    .X(_10362_));
 sky130_fd_sc_hd__nand2_1 _17344_ (.A(_10361_),
    .B(_10362_),
    .Y(_10363_));
 sky130_fd_sc_hd__a21oi_1 _17345_ (.A1(_10146_),
    .A2(_10238_),
    .B1(_10236_),
    .Y(_10364_));
 sky130_fd_sc_hd__xor2_1 _17346_ (.A(_10363_),
    .B(_10364_),
    .X(_10365_));
 sky130_fd_sc_hd__nand2_1 _17347_ (.A(_10144_),
    .B(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__or2_1 _17348_ (.A(_10144_),
    .B(_10365_),
    .X(_10367_));
 sky130_fd_sc_hd__nand2_1 _17349_ (.A(_10366_),
    .B(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__a21o_1 _17350_ (.A1(_10265_),
    .A2(_10242_),
    .B1(_10368_),
    .X(_10369_));
 sky130_fd_sc_hd__and3_1 _17351_ (.A(_10265_),
    .B(_10242_),
    .C(_10368_),
    .X(_10370_));
 sky130_fd_sc_hd__inv_2 _17352_ (.A(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__nand2_1 _17353_ (.A(_10369_),
    .B(_10371_),
    .Y(_10372_));
 sky130_fd_sc_hd__a21oi_1 _17354_ (.A1(_10246_),
    .A2(_10254_),
    .B1(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__a31o_1 _17355_ (.A1(_10246_),
    .A2(_10254_),
    .A3(_10372_),
    .B1(_08123_),
    .X(_10374_));
 sky130_fd_sc_hd__or2_2 _17356_ (.A(_10373_),
    .B(_10374_),
    .X(_10375_));
 sky130_fd_sc_hd__o311a_1 _17357_ (.A1(_09822_),
    .A2(_10263_),
    .A3(_10264_),
    .B1(_09812_),
    .C1(_10375_),
    .X(_10376_));
 sky130_fd_sc_hd__a21oi_1 _17358_ (.A1(_06171_),
    .A2(_09785_),
    .B1(_10376_),
    .Y(_00542_));
 sky130_fd_sc_hd__nand2_1 _17359_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .Y(_10377_));
 sky130_fd_sc_hd__or2_1 _17360_ (.A(\rbzero.wall_tracer.trackDistX[4] ),
    .B(\rbzero.wall_tracer.stepDistX[4] ),
    .X(_10378_));
 sky130_fd_sc_hd__o211a_1 _17361_ (.A1(_10261_),
    .A2(_10264_),
    .B1(_10377_),
    .C1(_10378_),
    .X(_10379_));
 sky130_fd_sc_hd__a211oi_1 _17362_ (.A1(_10377_),
    .A2(_10378_),
    .B1(_10261_),
    .C1(_10264_),
    .Y(_10380_));
 sky130_fd_sc_hd__or2b_1 _17363_ (.A(_10307_),
    .B_N(_10272_),
    .X(_10381_));
 sky130_fd_sc_hd__o2bb2a_1 _17364_ (.A1_N(_10284_),
    .A2_N(_10285_),
    .B1(_10282_),
    .B2(_10283_),
    .X(_10382_));
 sky130_fd_sc_hd__a21oi_2 _17365_ (.A1(_10305_),
    .A2(_10381_),
    .B1(_10382_),
    .Y(_10383_));
 sky130_fd_sc_hd__and3_1 _17366_ (.A(_10305_),
    .B(_10381_),
    .C(_10382_),
    .X(_10384_));
 sky130_fd_sc_hd__nor2_1 _17367_ (.A(_10383_),
    .B(_10384_),
    .Y(_10385_));
 sky130_fd_sc_hd__a21o_1 _17368_ (.A1(_10286_),
    .A2(_10303_),
    .B1(_10301_),
    .X(_10386_));
 sky130_fd_sc_hd__or2_1 _17369_ (.A(_10311_),
    .B(_10326_),
    .X(_10387_));
 sky130_fd_sc_hd__or2b_1 _17370_ (.A(_10327_),
    .B_N(_10309_),
    .X(_01663_));
 sky130_fd_sc_hd__nor2_1 _17371_ (.A(_09519_),
    .B(_09242_),
    .Y(_01664_));
 sky130_fd_sc_hd__xnor2_1 _17372_ (.A(_10275_),
    .B(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__or3_1 _17373_ (.A(_09525_),
    .B(_09491_),
    .C(_01665_),
    .X(_01666_));
 sky130_fd_sc_hd__o21ai_1 _17374_ (.A1(_09525_),
    .A2(_09491_),
    .B1(_01665_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _17375_ (.A(_01666_),
    .B(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__a21oi_1 _17376_ (.A1(_10150_),
    .A2(_10275_),
    .B1(_10280_),
    .Y(_01669_));
 sky130_fd_sc_hd__xor2_1 _17377_ (.A(_01668_),
    .B(_01669_),
    .X(_01670_));
 sky130_fd_sc_hd__and2_1 _17378_ (.A(_09146_),
    .B(_09687_),
    .X(_01671_));
 sky130_fd_sc_hd__xor2_1 _17379_ (.A(_01670_),
    .B(_01671_),
    .X(_01672_));
 sky130_fd_sc_hd__a21bo_1 _17380_ (.A1(_10291_),
    .A2(_10294_),
    .B1_N(_10292_),
    .X(_01673_));
 sky130_fd_sc_hd__or2b_1 _17381_ (.A(_10289_),
    .B_N(_10312_),
    .X(_01674_));
 sky130_fd_sc_hd__nand2_1 _17382_ (.A(_01674_),
    .B(_10314_),
    .Y(_01675_));
 sky130_fd_sc_hd__or2_1 _17383_ (.A(_08404_),
    .B(_09076_),
    .X(_01676_));
 sky130_fd_sc_hd__or3_1 _17384_ (.A(_08399_),
    .B(_08618_),
    .C(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__o21ai_1 _17385_ (.A1(_08399_),
    .A2(_08618_),
    .B1(_01676_),
    .Y(_01678_));
 sky130_fd_sc_hd__nand2_1 _17386_ (.A(_01677_),
    .B(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hd__nor2_1 _17387_ (.A(_09647_),
    .B(_09252_),
    .Y(_01680_));
 sky130_fd_sc_hd__xor2_1 _17388_ (.A(_01679_),
    .B(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__xnor2_1 _17389_ (.A(_01675_),
    .B(_01681_),
    .Y(_01682_));
 sky130_fd_sc_hd__xnor2_1 _17390_ (.A(_01673_),
    .B(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__a21oi_1 _17391_ (.A1(_10287_),
    .A2(_10298_),
    .B1(_10296_),
    .Y(_01684_));
 sky130_fd_sc_hd__nor2_1 _17392_ (.A(_01683_),
    .B(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__and2_1 _17393_ (.A(_01683_),
    .B(_01684_),
    .X(_01686_));
 sky130_fd_sc_hd__nor2_1 _17394_ (.A(_01685_),
    .B(_01686_),
    .Y(_01687_));
 sky130_fd_sc_hd__xnor2_1 _17395_ (.A(_01672_),
    .B(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__a21o_1 _17396_ (.A1(_10387_),
    .A2(_01663_),
    .B1(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__nand3_1 _17397_ (.A(_10387_),
    .B(_01663_),
    .C(_01688_),
    .Y(_01690_));
 sky130_fd_sc_hd__nand2_1 _17398_ (.A(_01689_),
    .B(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__xnor2_1 _17399_ (.A(_10386_),
    .B(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__nor2_1 _17400_ (.A(_10322_),
    .B(_10324_),
    .Y(_01693_));
 sky130_fd_sc_hd__a21o_1 _17401_ (.A1(_10317_),
    .A2(_10325_),
    .B1(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__or2b_1 _17402_ (.A(_10338_),
    .B_N(_10329_),
    .X(_01695_));
 sky130_fd_sc_hd__a21bo_1 _17403_ (.A1(_10332_),
    .A2(_10337_),
    .B1_N(_01695_),
    .X(_01696_));
 sky130_fd_sc_hd__nand2_2 _17404_ (.A(\rbzero.wall_tracer.visualWallDist[1] ),
    .B(_08421_),
    .Y(_01697_));
 sky130_fd_sc_hd__or4_1 _17405_ (.A(_01697_),
    .B(_10288_),
    .C(_08476_),
    .D(_09044_),
    .X(_01698_));
 sky130_fd_sc_hd__and2_1 _17406_ (.A(_08475_),
    .B(_08445_),
    .X(_01699_));
 sky130_fd_sc_hd__nor2_1 _17407_ (.A(_01697_),
    .B(_09044_),
    .Y(_01700_));
 sky130_fd_sc_hd__a31o_1 _17408_ (.A1(\rbzero.wall_tracer.visualWallDist[2] ),
    .A2(_08421_),
    .A3(_01699_),
    .B1(_01700_),
    .X(_01701_));
 sky130_fd_sc_hd__nand2_1 _17409_ (.A(_01698_),
    .B(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__or2_1 _17410_ (.A(_08499_),
    .B(_08620_),
    .X(_01703_));
 sky130_fd_sc_hd__xor2_2 _17411_ (.A(_01702_),
    .B(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__nor2_1 _17412_ (.A(_08814_),
    .B(_09677_),
    .Y(_01705_));
 sky130_fd_sc_hd__xnor2_1 _17413_ (.A(_10318_),
    .B(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__nor2_1 _17414_ (.A(_09397_),
    .B(_09186_),
    .Y(_01707_));
 sky130_fd_sc_hd__xor2_1 _17415_ (.A(_01706_),
    .B(_01707_),
    .X(_01708_));
 sky130_fd_sc_hd__a22oi_2 _17416_ (.A1(_10190_),
    .A2(_10318_),
    .B1(_10320_),
    .B2(_10321_),
    .Y(_01709_));
 sky130_fd_sc_hd__xor2_1 _17417_ (.A(_01708_),
    .B(_01709_),
    .X(_01710_));
 sky130_fd_sc_hd__nand2_1 _17418_ (.A(_01704_),
    .B(_01710_),
    .Y(_01711_));
 sky130_fd_sc_hd__or2_1 _17419_ (.A(_01704_),
    .B(_01710_),
    .X(_01712_));
 sky130_fd_sc_hd__nand2_1 _17420_ (.A(_01711_),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__xor2_1 _17421_ (.A(_01696_),
    .B(_01713_),
    .X(_01714_));
 sky130_fd_sc_hd__xnor2_1 _17422_ (.A(_01694_),
    .B(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hd__or3_1 _17423_ (.A(_09542_),
    .B(_09677_),
    .C(_10335_),
    .X(_01716_));
 sky130_fd_sc_hd__a21bo_1 _17424_ (.A1(_10333_),
    .A2(_10334_),
    .B1_N(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__buf_2 _17425_ (.A(_10330_),
    .X(_01718_));
 sky130_fd_sc_hd__o31ai_1 _17426_ (.A1(_09167_),
    .A2(_01718_),
    .A3(_10342_),
    .B1(_10331_),
    .Y(_01719_));
 sky130_fd_sc_hd__or2_1 _17427_ (.A(_08816_),
    .B(_10215_),
    .X(_01720_));
 sky130_fd_sc_hd__nor2_1 _17428_ (.A(_08889_),
    .B(_10330_),
    .Y(_01721_));
 sky130_fd_sc_hd__xor2_1 _17429_ (.A(_01720_),
    .B(_01721_),
    .X(_01722_));
 sky130_fd_sc_hd__nor2_1 _17430_ (.A(_09542_),
    .B(_09560_),
    .Y(_01723_));
 sky130_fd_sc_hd__xor2_1 _17431_ (.A(_01722_),
    .B(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__xor2_1 _17432_ (.A(_01719_),
    .B(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__xnor2_1 _17433_ (.A(_01717_),
    .B(_01725_),
    .Y(_01726_));
 sky130_fd_sc_hd__a21o_1 _17434_ (.A1(_10096_),
    .A2(_10344_),
    .B1(_10221_),
    .X(_01727_));
 sky130_fd_sc_hd__nor2_1 _17435_ (.A(_09167_),
    .B(_10093_),
    .Y(_01728_));
 sky130_fd_sc_hd__mux2_2 _17436_ (.A0(_09167_),
    .A1(_01728_),
    .S(_10342_),
    .X(_01729_));
 sky130_fd_sc_hd__xor2_1 _17437_ (.A(_10096_),
    .B(_01729_),
    .X(_01730_));
 sky130_fd_sc_hd__and2_1 _17438_ (.A(_01727_),
    .B(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__nor2_1 _17439_ (.A(_01727_),
    .B(_01730_),
    .Y(_01732_));
 sky130_fd_sc_hd__nor2_1 _17440_ (.A(_01731_),
    .B(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__xnor2_1 _17441_ (.A(_01726_),
    .B(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__nor2_1 _17442_ (.A(_10345_),
    .B(_10346_),
    .Y(_01735_));
 sky130_fd_sc_hd__a21oi_1 _17443_ (.A1(_10339_),
    .A2(_10347_),
    .B1(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__xor2_1 _17444_ (.A(_01734_),
    .B(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__xnor2_1 _17445_ (.A(_01715_),
    .B(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__and2b_1 _17446_ (.A_N(_10348_),
    .B(_10350_),
    .X(_01739_));
 sky130_fd_sc_hd__a21oi_1 _17447_ (.A1(_10328_),
    .A2(_10351_),
    .B1(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__xor2_1 _17448_ (.A(_01738_),
    .B(_01740_),
    .X(_01741_));
 sky130_fd_sc_hd__xnor2_1 _17449_ (.A(_01692_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__a21oi_1 _17450_ (.A1(_10308_),
    .A2(_10357_),
    .B1(_10355_),
    .Y(_01743_));
 sky130_fd_sc_hd__nor2_1 _17451_ (.A(_01742_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__nand2_1 _17452_ (.A(_01742_),
    .B(_01743_),
    .Y(_01745_));
 sky130_fd_sc_hd__and2b_1 _17453_ (.A_N(_01744_),
    .B(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__xnor2_1 _17454_ (.A(_10385_),
    .B(_01746_),
    .Y(_01747_));
 sky130_fd_sc_hd__o21a_1 _17455_ (.A1(_10358_),
    .A2(_10359_),
    .B1(_10361_),
    .X(_01748_));
 sky130_fd_sc_hd__xor2_1 _17456_ (.A(_01747_),
    .B(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__nand2_1 _17457_ (.A(_10269_),
    .B(_01749_),
    .Y(_01750_));
 sky130_fd_sc_hd__or2_1 _17458_ (.A(_10269_),
    .B(_01749_),
    .X(_01751_));
 sky130_fd_sc_hd__nand2_2 _17459_ (.A(_01750_),
    .B(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hd__o21a_1 _17460_ (.A1(_10363_),
    .A2(_10364_),
    .B1(_10366_),
    .X(_01753_));
 sky130_fd_sc_hd__xor2_4 _17461_ (.A(_01752_),
    .B(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__a21oi_1 _17462_ (.A1(_10246_),
    .A2(_10369_),
    .B1(_10370_),
    .Y(_01755_));
 sky130_fd_sc_hd__a41o_1 _17463_ (.A1(_10248_),
    .A2(_10253_),
    .A3(_10369_),
    .A4(_10371_),
    .B1(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__buf_8 _17464_ (.A(_08123_),
    .X(_01757_));
 sky130_fd_sc_hd__a21oi_1 _17465_ (.A1(_01754_),
    .A2(_01756_),
    .B1(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__o21ai_4 _17466_ (.A1(_01754_),
    .A2(_01756_),
    .B1(_01758_),
    .Y(_01759_));
 sky130_fd_sc_hd__o311a_1 _17467_ (.A1(_09822_),
    .A2(_10379_),
    .A3(_10380_),
    .B1(_09812_),
    .C1(_01759_),
    .X(_01760_));
 sky130_fd_sc_hd__a21oi_1 _17468_ (.A1(_06170_),
    .A2(_09785_),
    .B1(_01760_),
    .Y(_00543_));
 sky130_fd_sc_hd__nor2_1 _17469_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .Y(_01761_));
 sky130_fd_sc_hd__and2_1 _17470_ (.A(\rbzero.wall_tracer.trackDistX[5] ),
    .B(\rbzero.wall_tracer.stepDistX[5] ),
    .X(_01762_));
 sky130_fd_sc_hd__a21oi_1 _17471_ (.A1(\rbzero.wall_tracer.trackDistX[4] ),
    .A2(\rbzero.wall_tracer.stepDistX[4] ),
    .B1(_10379_),
    .Y(_01763_));
 sky130_fd_sc_hd__nor3_1 _17472_ (.A(_01761_),
    .B(_01762_),
    .C(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__o21a_1 _17473_ (.A1(_01761_),
    .A2(_01762_),
    .B1(_01763_),
    .X(_01765_));
 sky130_fd_sc_hd__or2_1 _17474_ (.A(_01747_),
    .B(_01748_),
    .X(_01766_));
 sky130_fd_sc_hd__or2b_1 _17475_ (.A(_01691_),
    .B_N(_10386_),
    .X(_01767_));
 sky130_fd_sc_hd__o2bb2a_1 _17476_ (.A1_N(_01670_),
    .A2_N(_01671_),
    .B1(_01668_),
    .B2(_01669_),
    .X(_01768_));
 sky130_fd_sc_hd__a21oi_1 _17477_ (.A1(_01689_),
    .A2(_01767_),
    .B1(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__and3_1 _17478_ (.A(_01689_),
    .B(_01767_),
    .C(_01768_),
    .X(_01770_));
 sky130_fd_sc_hd__nor2_1 _17479_ (.A(_01769_),
    .B(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__a21o_1 _17480_ (.A1(_01672_),
    .A2(_01687_),
    .B1(_01685_),
    .X(_01772_));
 sky130_fd_sc_hd__or2b_1 _17481_ (.A(_01713_),
    .B_N(_01696_),
    .X(_01773_));
 sky130_fd_sc_hd__or2b_1 _17482_ (.A(_01714_),
    .B_N(_01694_),
    .X(_01774_));
 sky130_fd_sc_hd__o22a_1 _17483_ (.A1(_09647_),
    .A2(_09243_),
    .B1(_09363_),
    .B2(_09519_),
    .X(_01775_));
 sky130_fd_sc_hd__or2_1 _17484_ (.A(_09647_),
    .B(_09362_),
    .X(_01776_));
 sky130_fd_sc_hd__or3_1 _17485_ (.A(_09519_),
    .B(_09242_),
    .C(_01776_),
    .X(_01777_));
 sky130_fd_sc_hd__and2b_1 _17486_ (.A_N(_01775_),
    .B(_01777_),
    .X(_01778_));
 sky130_fd_sc_hd__nor2_1 _17487_ (.A(_09520_),
    .B(_09491_),
    .Y(_01779_));
 sky130_fd_sc_hd__xnor2_1 _17488_ (.A(_01778_),
    .B(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__o31a_1 _17489_ (.A1(_09519_),
    .A2(_09363_),
    .A3(_10276_),
    .B1(_01666_),
    .X(_01781_));
 sky130_fd_sc_hd__xnor2_1 _17490_ (.A(_01780_),
    .B(_01781_),
    .Y(_01782_));
 sky130_fd_sc_hd__nand2_1 _17491_ (.A(_09525_),
    .B(_09890_),
    .Y(_01783_));
 sky130_fd_sc_hd__xor2_1 _17492_ (.A(_01782_),
    .B(_01783_),
    .X(_01784_));
 sky130_fd_sc_hd__o31ai_2 _17493_ (.A1(_09647_),
    .A2(_09252_),
    .A3(_01679_),
    .B1(_01677_),
    .Y(_01785_));
 sky130_fd_sc_hd__o21ai_1 _17494_ (.A1(_01702_),
    .A2(_01703_),
    .B1(_01698_),
    .Y(_01786_));
 sky130_fd_sc_hd__or2_1 _17495_ (.A(_08499_),
    .B(_08617_),
    .X(_01787_));
 sky130_fd_sc_hd__or3_1 _17496_ (.A(_08399_),
    .B(_09079_),
    .C(_01787_),
    .X(_01788_));
 sky130_fd_sc_hd__o21ai_1 _17497_ (.A1(_10315_),
    .A2(_09079_),
    .B1(_01787_),
    .Y(_01789_));
 sky130_fd_sc_hd__nand2_1 _17498_ (.A(_01788_),
    .B(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__nor2_1 _17499_ (.A(_10059_),
    .B(_09252_),
    .Y(_01791_));
 sky130_fd_sc_hd__xor2_1 _17500_ (.A(_01790_),
    .B(_01791_),
    .X(_01792_));
 sky130_fd_sc_hd__xnor2_1 _17501_ (.A(_01786_),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__xnor2_1 _17502_ (.A(_01785_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__a21oi_1 _17503_ (.A1(_01674_),
    .A2(_10314_),
    .B1(_01681_),
    .Y(_01795_));
 sky130_fd_sc_hd__a21oi_1 _17504_ (.A1(_01673_),
    .A2(_01682_),
    .B1(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__nor2_1 _17505_ (.A(_01794_),
    .B(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__and2_1 _17506_ (.A(_01794_),
    .B(_01796_),
    .X(_01798_));
 sky130_fd_sc_hd__nor2_1 _17507_ (.A(_01797_),
    .B(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__xnor2_1 _17508_ (.A(_01784_),
    .B(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__a21o_1 _17509_ (.A1(_01773_),
    .A2(_01774_),
    .B1(_01800_),
    .X(_01801_));
 sky130_fd_sc_hd__nand3_1 _17510_ (.A(_01773_),
    .B(_01774_),
    .C(_01800_),
    .Y(_01802_));
 sky130_fd_sc_hd__nand2_1 _17511_ (.A(_01801_),
    .B(_01802_),
    .Y(_01803_));
 sky130_fd_sc_hd__xnor2_1 _17512_ (.A(_01772_),
    .B(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__o21ai_1 _17513_ (.A1(_01708_),
    .A2(_01709_),
    .B1(_01711_),
    .Y(_01805_));
 sky130_fd_sc_hd__or2b_1 _17514_ (.A(_01724_),
    .B_N(_01719_),
    .X(_01806_));
 sky130_fd_sc_hd__or2b_1 _17515_ (.A(_01725_),
    .B_N(_01717_),
    .X(_01807_));
 sky130_fd_sc_hd__nand2_1 _17516_ (.A(_01806_),
    .B(_01807_),
    .Y(_01808_));
 sky130_fd_sc_hd__nor2_2 _17517_ (.A(_10288_),
    .B(_09670_),
    .Y(_01809_));
 sky130_fd_sc_hd__o22a_1 _17518_ (.A1(_10288_),
    .A2(_09662_),
    .B1(_09670_),
    .B2(_01697_),
    .X(_01810_));
 sky130_fd_sc_hd__a21oi_2 _17519_ (.A1(_01700_),
    .A2(_01809_),
    .B1(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__and3_1 _17520_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08475_),
    .C(_08445_),
    .X(_01812_));
 sky130_fd_sc_hd__xor2_2 _17521_ (.A(_01811_),
    .B(_01812_),
    .X(_01813_));
 sky130_fd_sc_hd__or2_1 _17522_ (.A(_09528_),
    .B(_09559_),
    .X(_01814_));
 sky130_fd_sc_hd__or3_1 _17523_ (.A(_08814_),
    .B(_09677_),
    .C(_01814_),
    .X(_01815_));
 sky130_fd_sc_hd__o22ai_1 _17524_ (.A1(_09528_),
    .A2(_09677_),
    .B1(_09560_),
    .B2(_08814_),
    .Y(_01816_));
 sky130_fd_sc_hd__nand2_1 _17525_ (.A(_01815_),
    .B(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__buf_2 _17526_ (.A(_09397_),
    .X(_01818_));
 sky130_fd_sc_hd__nor2_1 _17527_ (.A(_01818_),
    .B(_09669_),
    .Y(_01819_));
 sky130_fd_sc_hd__xor2_1 _17528_ (.A(_01817_),
    .B(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__nand2_1 _17529_ (.A(_10318_),
    .B(_01705_),
    .Y(_01821_));
 sky130_fd_sc_hd__o31a_1 _17530_ (.A1(_01818_),
    .A2(_09186_),
    .A3(_01706_),
    .B1(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__nor2_1 _17531_ (.A(_01820_),
    .B(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__and2_1 _17532_ (.A(_01820_),
    .B(_01822_),
    .X(_01824_));
 sky130_fd_sc_hd__nor2_1 _17533_ (.A(_01823_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__xnor2_1 _17534_ (.A(_01813_),
    .B(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__xor2_1 _17535_ (.A(_01808_),
    .B(_01826_),
    .X(_01827_));
 sky130_fd_sc_hd__xnor2_1 _17536_ (.A(_01805_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__or3_1 _17537_ (.A(_08889_),
    .B(_01718_),
    .C(_01720_),
    .X(_01829_));
 sky130_fd_sc_hd__o31ai_1 _17538_ (.A1(_09542_),
    .A2(_09560_),
    .A3(_01722_),
    .B1(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__o21ai_4 _17539_ (.A1(_09167_),
    .A2(_10342_),
    .B1(_10331_),
    .Y(_01831_));
 sky130_fd_sc_hd__or3_2 _17540_ (.A(_08889_),
    .B(_08816_),
    .C(_10093_),
    .X(_01832_));
 sky130_fd_sc_hd__o22ai_1 _17541_ (.A1(_08889_),
    .A2(_10093_),
    .B1(_10330_),
    .B2(_08816_),
    .Y(_01833_));
 sky130_fd_sc_hd__o21ai_1 _17542_ (.A1(_01718_),
    .A2(_01832_),
    .B1(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__nor2_1 _17543_ (.A(_09542_),
    .B(_10215_),
    .Y(_01835_));
 sky130_fd_sc_hd__xnor2_1 _17544_ (.A(_01834_),
    .B(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__xnor2_1 _17545_ (.A(_01831_),
    .B(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__xnor2_1 _17546_ (.A(_01830_),
    .B(_01837_),
    .Y(_01838_));
 sky130_fd_sc_hd__nand2_1 _17547_ (.A(_10221_),
    .B(_01729_),
    .Y(_01839_));
 sky130_fd_sc_hd__or2_1 _17548_ (.A(_10094_),
    .B(_01729_),
    .X(_01840_));
 sky130_fd_sc_hd__and2_1 _17549_ (.A(_01839_),
    .B(_01840_),
    .X(_01841_));
 sky130_fd_sc_hd__buf_2 _17550_ (.A(_01841_),
    .X(_01842_));
 sky130_fd_sc_hd__xnor2_1 _17551_ (.A(_01838_),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__a21oi_1 _17552_ (.A1(_01726_),
    .A2(_01733_),
    .B1(_01731_),
    .Y(_01844_));
 sky130_fd_sc_hd__nor2_1 _17553_ (.A(_01843_),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__and2_1 _17554_ (.A(_01843_),
    .B(_01844_),
    .X(_01846_));
 sky130_fd_sc_hd__nor2_1 _17555_ (.A(_01845_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__xnor2_1 _17556_ (.A(_01828_),
    .B(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor2_1 _17557_ (.A(_01734_),
    .B(_01736_),
    .Y(_01849_));
 sky130_fd_sc_hd__a21oi_1 _17558_ (.A1(_01715_),
    .A2(_01737_),
    .B1(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__xor2_1 _17559_ (.A(_01848_),
    .B(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__xnor2_1 _17560_ (.A(_01804_),
    .B(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__nor2_1 _17561_ (.A(_01738_),
    .B(_01740_),
    .Y(_01853_));
 sky130_fd_sc_hd__a21oi_1 _17562_ (.A1(_01692_),
    .A2(_01741_),
    .B1(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__xor2_1 _17563_ (.A(_01852_),
    .B(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__xnor2_1 _17564_ (.A(_01771_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__a21oi_1 _17565_ (.A1(_10385_),
    .A2(_01745_),
    .B1(_01744_),
    .Y(_01857_));
 sky130_fd_sc_hd__nor2_1 _17566_ (.A(_01856_),
    .B(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand2_1 _17567_ (.A(_01856_),
    .B(_01857_),
    .Y(_01859_));
 sky130_fd_sc_hd__and2b_1 _17568_ (.A_N(_01858_),
    .B(_01859_),
    .X(_01860_));
 sky130_fd_sc_hd__xnor2_1 _17569_ (.A(_10383_),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__and3_1 _17570_ (.A(_01766_),
    .B(_01750_),
    .C(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__a21oi_1 _17571_ (.A1(_01766_),
    .A2(_01750_),
    .B1(_01861_),
    .Y(_01863_));
 sky130_fd_sc_hd__or2_1 _17572_ (.A(_01862_),
    .B(_01863_),
    .X(_01864_));
 sky130_fd_sc_hd__or2_1 _17573_ (.A(_01752_),
    .B(_01753_),
    .X(_01865_));
 sky130_fd_sc_hd__a21boi_2 _17574_ (.A1(_01754_),
    .A2(_01756_),
    .B1_N(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__a21oi_1 _17575_ (.A1(_01864_),
    .A2(_01866_),
    .B1(_01757_),
    .Y(_01867_));
 sky130_fd_sc_hd__o21ai_4 _17576_ (.A1(_01864_),
    .A2(_01866_),
    .B1(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__o311a_1 _17577_ (.A1(_09822_),
    .A2(_01764_),
    .A3(_01765_),
    .B1(_09812_),
    .C1(_01868_),
    .X(_01869_));
 sky130_fd_sc_hd__a21oi_1 _17578_ (.A1(_06169_),
    .A2(_09785_),
    .B1(_01869_),
    .Y(_00544_));
 sky130_fd_sc_hd__nor2_1 _17579_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_01870_));
 sky130_fd_sc_hd__nand2_1 _17580_ (.A(\rbzero.wall_tracer.trackDistX[6] ),
    .B(\rbzero.wall_tracer.stepDistX[6] ),
    .Y(_01871_));
 sky130_fd_sc_hd__or2b_1 _17581_ (.A(_01870_),
    .B_N(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__o21ba_1 _17582_ (.A1(_01761_),
    .A2(_01763_),
    .B1_N(_01762_),
    .X(_01873_));
 sky130_fd_sc_hd__nor2_1 _17583_ (.A(_01872_),
    .B(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__a21o_1 _17584_ (.A1(_01872_),
    .A2(_01873_),
    .B1(_09866_),
    .X(_01875_));
 sky130_fd_sc_hd__or2b_1 _17585_ (.A(_01803_),
    .B_N(_01772_),
    .X(_01876_));
 sky130_fd_sc_hd__o22a_1 _17586_ (.A1(_01780_),
    .A2(_01781_),
    .B1(_01782_),
    .B2(_01783_),
    .X(_01877_));
 sky130_fd_sc_hd__a21oi_2 _17587_ (.A1(_01801_),
    .A2(_01876_),
    .B1(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__and3_1 _17588_ (.A(_01801_),
    .B(_01876_),
    .C(_01877_),
    .X(_01879_));
 sky130_fd_sc_hd__nor2_1 _17589_ (.A(_01878_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__a21o_1 _17590_ (.A1(_01784_),
    .A2(_01799_),
    .B1(_01797_),
    .X(_01881_));
 sky130_fd_sc_hd__or2b_1 _17591_ (.A(_01826_),
    .B_N(_01808_),
    .X(_01882_));
 sky130_fd_sc_hd__or2b_1 _17592_ (.A(_01827_),
    .B_N(_01805_),
    .X(_01883_));
 sky130_fd_sc_hd__nor2_1 _17593_ (.A(_10059_),
    .B(_09243_),
    .Y(_01884_));
 sky130_fd_sc_hd__xnor2_1 _17594_ (.A(_01776_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__nor2_1 _17595_ (.A(_09519_),
    .B(_09621_),
    .Y(_01886_));
 sky130_fd_sc_hd__nand2_1 _17596_ (.A(_01885_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__or2_1 _17597_ (.A(_01885_),
    .B(_01886_),
    .X(_01888_));
 sky130_fd_sc_hd__nand2_1 _17598_ (.A(_01887_),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__o31a_1 _17599_ (.A1(_09520_),
    .A2(_09621_),
    .A3(_01775_),
    .B1(_01777_),
    .X(_01890_));
 sky130_fd_sc_hd__xor2_2 _17600_ (.A(_01889_),
    .B(_01890_),
    .X(_01891_));
 sky130_fd_sc_hd__and2_1 _17601_ (.A(_09520_),
    .B(_09890_),
    .X(_01892_));
 sky130_fd_sc_hd__xor2_2 _17602_ (.A(_01891_),
    .B(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__o31ai_2 _17603_ (.A1(_10059_),
    .A2(_09252_),
    .A3(_01790_),
    .B1(_01788_),
    .Y(_01894_));
 sky130_fd_sc_hd__nand2_1 _17604_ (.A(_01700_),
    .B(_01809_),
    .Y(_01895_));
 sky130_fd_sc_hd__nand2_1 _17605_ (.A(_01811_),
    .B(_01812_),
    .Y(_01896_));
 sky130_fd_sc_hd__or2_1 _17606_ (.A(_10315_),
    .B(_09252_),
    .X(_01897_));
 sky130_fd_sc_hd__nand2_1 _17607_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_08421_),
    .Y(_01898_));
 sky130_fd_sc_hd__nor2_1 _17608_ (.A(_08428_),
    .B(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__a31o_1 _17609_ (.A1(\rbzero.wall_tracer.visualWallDist[4] ),
    .A2(_08421_),
    .A3(_01699_),
    .B1(_01899_),
    .X(_01900_));
 sky130_fd_sc_hd__nand2_1 _17610_ (.A(\rbzero.wall_tracer.visualWallDist[5] ),
    .B(_01699_),
    .Y(_01901_));
 sky130_fd_sc_hd__or2_1 _17611_ (.A(_01787_),
    .B(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__nand2_1 _17612_ (.A(_01900_),
    .B(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__xnor2_1 _17613_ (.A(_01897_),
    .B(_01903_),
    .Y(_01904_));
 sky130_fd_sc_hd__a21oi_1 _17614_ (.A1(_01895_),
    .A2(_01896_),
    .B1(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__and3_1 _17615_ (.A(_01895_),
    .B(_01896_),
    .C(_01904_),
    .X(_01906_));
 sky130_fd_sc_hd__nor2_1 _17616_ (.A(_01905_),
    .B(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__xnor2_1 _17617_ (.A(_01894_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__and2b_1 _17618_ (.A_N(_01792_),
    .B(_01786_),
    .X(_01909_));
 sky130_fd_sc_hd__a21oi_1 _17619_ (.A1(_01785_),
    .A2(_01793_),
    .B1(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__nor2_1 _17620_ (.A(_01908_),
    .B(_01910_),
    .Y(_01911_));
 sky130_fd_sc_hd__and2_1 _17621_ (.A(_01908_),
    .B(_01910_),
    .X(_01912_));
 sky130_fd_sc_hd__nor2_1 _17622_ (.A(_01911_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__xnor2_2 _17623_ (.A(_01893_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__a21o_1 _17624_ (.A1(_01882_),
    .A2(_01883_),
    .B1(_01914_),
    .X(_01915_));
 sky130_fd_sc_hd__nand3_1 _17625_ (.A(_01882_),
    .B(_01883_),
    .C(_01914_),
    .Y(_01916_));
 sky130_fd_sc_hd__nand2_1 _17626_ (.A(_01915_),
    .B(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__xnor2_1 _17627_ (.A(_01881_),
    .B(_01917_),
    .Y(_01918_));
 sky130_fd_sc_hd__a21o_1 _17628_ (.A1(_01813_),
    .A2(_01825_),
    .B1(_01823_),
    .X(_01919_));
 sky130_fd_sc_hd__nand2_1 _17629_ (.A(_01831_),
    .B(_01836_),
    .Y(_01920_));
 sky130_fd_sc_hd__or2b_1 _17630_ (.A(_01837_),
    .B_N(_01830_),
    .X(_01921_));
 sky130_fd_sc_hd__nand2_2 _17631_ (.A(\rbzero.wall_tracer.visualWallDist[3] ),
    .B(_08421_),
    .Y(_01922_));
 sky130_fd_sc_hd__nor2_1 _17632_ (.A(_01697_),
    .B(_09315_),
    .Y(_01923_));
 sky130_fd_sc_hd__xnor2_1 _17633_ (.A(_01809_),
    .B(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__or3_1 _17634_ (.A(_09662_),
    .B(_01922_),
    .C(_01924_),
    .X(_01925_));
 sky130_fd_sc_hd__o21ai_1 _17635_ (.A1(_09662_),
    .A2(_01922_),
    .B1(_01924_),
    .Y(_01926_));
 sky130_fd_sc_hd__and2_1 _17636_ (.A(_01925_),
    .B(_01926_),
    .X(_01927_));
 sky130_fd_sc_hd__or2_1 _17637_ (.A(_08814_),
    .B(_10215_),
    .X(_01928_));
 sky130_fd_sc_hd__xnor2_1 _17638_ (.A(_01814_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__nor2_1 _17639_ (.A(_01818_),
    .B(_09677_),
    .Y(_01930_));
 sky130_fd_sc_hd__xor2_1 _17640_ (.A(_01929_),
    .B(_01930_),
    .X(_01931_));
 sky130_fd_sc_hd__o31a_1 _17641_ (.A1(_01818_),
    .A2(_09669_),
    .A3(_01817_),
    .B1(_01815_),
    .X(_01932_));
 sky130_fd_sc_hd__nor2_1 _17642_ (.A(_01931_),
    .B(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__and2_1 _17643_ (.A(_01931_),
    .B(_01932_),
    .X(_01934_));
 sky130_fd_sc_hd__nor2_1 _17644_ (.A(_01933_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__xnor2_1 _17645_ (.A(_01927_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__a21o_1 _17646_ (.A1(_01920_),
    .A2(_01921_),
    .B1(_01936_),
    .X(_01937_));
 sky130_fd_sc_hd__nand3_1 _17647_ (.A(_01920_),
    .B(_01921_),
    .C(_01936_),
    .Y(_01938_));
 sky130_fd_sc_hd__nand2_1 _17648_ (.A(_01937_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__xnor2_1 _17649_ (.A(_01919_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__a2bb2o_1 _17650_ (.A1_N(_01718_),
    .A2_N(_01832_),
    .B1(_01835_),
    .B2(_01833_),
    .X(_01941_));
 sky130_fd_sc_hd__and2_1 _17651_ (.A(_08889_),
    .B(_08816_),
    .X(_01942_));
 sky130_fd_sc_hd__or3b_1 _17652_ (.A(_01942_),
    .B(_10093_),
    .C_N(_01832_),
    .X(_01943_));
 sky130_fd_sc_hd__nor2_1 _17653_ (.A(_09542_),
    .B(_01718_),
    .Y(_01944_));
 sky130_fd_sc_hd__xnor2_1 _17654_ (.A(_01943_),
    .B(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__and2_1 _17655_ (.A(_01831_),
    .B(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__nor2_1 _17656_ (.A(_01831_),
    .B(_01945_),
    .Y(_01947_));
 sky130_fd_sc_hd__nor2_1 _17657_ (.A(_01946_),
    .B(_01947_),
    .Y(_01948_));
 sky130_fd_sc_hd__xor2_1 _17658_ (.A(_01941_),
    .B(_01948_),
    .X(_01949_));
 sky130_fd_sc_hd__xnor2_1 _17659_ (.A(_01842_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__a21boi_1 _17660_ (.A1(_01838_),
    .A2(_01842_),
    .B1_N(_01839_),
    .Y(_01951_));
 sky130_fd_sc_hd__nor2_1 _17661_ (.A(_01950_),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__and2_1 _17662_ (.A(_01950_),
    .B(_01951_),
    .X(_01953_));
 sky130_fd_sc_hd__nor2_1 _17663_ (.A(_01952_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__xnor2_1 _17664_ (.A(_01940_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__a21oi_1 _17665_ (.A1(_01828_),
    .A2(_01847_),
    .B1(_01845_),
    .Y(_01956_));
 sky130_fd_sc_hd__xor2_1 _17666_ (.A(_01955_),
    .B(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__xnor2_1 _17667_ (.A(_01918_),
    .B(_01957_),
    .Y(_01958_));
 sky130_fd_sc_hd__nor2_1 _17668_ (.A(_01848_),
    .B(_01850_),
    .Y(_01959_));
 sky130_fd_sc_hd__a21oi_1 _17669_ (.A1(_01804_),
    .A2(_01851_),
    .B1(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__xor2_1 _17670_ (.A(_01958_),
    .B(_01960_),
    .X(_01961_));
 sky130_fd_sc_hd__xnor2_1 _17671_ (.A(_01880_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_1 _17672_ (.A(_01852_),
    .B(_01854_),
    .Y(_01963_));
 sky130_fd_sc_hd__a21oi_1 _17673_ (.A1(_01771_),
    .A2(_01855_),
    .B1(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__or2_1 _17674_ (.A(_01962_),
    .B(_01964_),
    .X(_01965_));
 sky130_fd_sc_hd__nand2_1 _17675_ (.A(_01962_),
    .B(_01964_),
    .Y(_01966_));
 sky130_fd_sc_hd__and2_1 _17676_ (.A(_01965_),
    .B(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__nand2_1 _17677_ (.A(_01769_),
    .B(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__or2_1 _17678_ (.A(_01769_),
    .B(_01967_),
    .X(_01969_));
 sky130_fd_sc_hd__nand2_1 _17679_ (.A(_01968_),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hd__a21oi_4 _17680_ (.A1(_10383_),
    .A2(_01859_),
    .B1(_01858_),
    .Y(_01971_));
 sky130_fd_sc_hd__or2_1 _17681_ (.A(_01970_),
    .B(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__nand2_1 _17682_ (.A(_01970_),
    .B(_01971_),
    .Y(_01973_));
 sky130_fd_sc_hd__nand2_1 _17683_ (.A(_01972_),
    .B(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__or3b_1 _17684_ (.A(_01862_),
    .B(_01863_),
    .C_N(_01754_),
    .X(_01975_));
 sky130_fd_sc_hd__or2b_1 _17685_ (.A(_01975_),
    .B_N(_01755_),
    .X(_01976_));
 sky130_fd_sc_hd__o41a_2 _17686_ (.A1(_10255_),
    .A2(_10256_),
    .A3(_10372_),
    .A4(_01975_),
    .B1(_01976_),
    .X(_01977_));
 sky130_fd_sc_hd__o21ba_2 _17687_ (.A1(_01865_),
    .A2(_01862_),
    .B1_N(_01863_),
    .X(_01978_));
 sky130_fd_sc_hd__and3_1 _17688_ (.A(_01974_),
    .B(_01977_),
    .C(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__a21o_1 _17689_ (.A1(_01977_),
    .A2(_01978_),
    .B1(_01974_),
    .X(_01980_));
 sky130_fd_sc_hd__or3b_1 _17690_ (.A(_08123_),
    .B(_01979_),
    .C_N(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__o21ai_1 _17691_ (.A1(_01874_),
    .A2(_01875_),
    .B1(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__mux2_1 _17692_ (.A0(\rbzero.wall_tracer.trackDistX[6] ),
    .A1(_01982_),
    .S(_09844_),
    .X(_01983_));
 sky130_fd_sc_hd__clkbuf_1 _17693_ (.A(_01983_),
    .X(_00545_));
 sky130_fd_sc_hd__nor2_1 _17694_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_01984_));
 sky130_fd_sc_hd__nand2_1 _17695_ (.A(\rbzero.wall_tracer.trackDistX[7] ),
    .B(\rbzero.wall_tracer.stepDistX[7] ),
    .Y(_01985_));
 sky130_fd_sc_hd__or2b_1 _17696_ (.A(_01984_),
    .B_N(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__o21a_1 _17697_ (.A1(_01870_),
    .A2(_01873_),
    .B1(_01871_),
    .X(_01987_));
 sky130_fd_sc_hd__nor2_1 _17698_ (.A(_01986_),
    .B(_01987_),
    .Y(_01988_));
 sky130_fd_sc_hd__a21o_1 _17699_ (.A1(_01986_),
    .A2(_01987_),
    .B1(_09866_),
    .X(_01989_));
 sky130_fd_sc_hd__or2b_1 _17700_ (.A(_01917_),
    .B_N(_01881_),
    .X(_01990_));
 sky130_fd_sc_hd__o2bb2a_1 _17701_ (.A1_N(_01891_),
    .A2_N(_01892_),
    .B1(_01889_),
    .B2(_01890_),
    .X(_01991_));
 sky130_fd_sc_hd__a21oi_2 _17702_ (.A1(_01915_),
    .A2(_01990_),
    .B1(_01991_),
    .Y(_01992_));
 sky130_fd_sc_hd__and3_1 _17703_ (.A(_01915_),
    .B(_01990_),
    .C(_01991_),
    .X(_01993_));
 sky130_fd_sc_hd__nor2_1 _17704_ (.A(_01992_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__a21o_1 _17705_ (.A1(_01893_),
    .A2(_01913_),
    .B1(_01911_),
    .X(_01995_));
 sky130_fd_sc_hd__or2b_1 _17706_ (.A(_01939_),
    .B_N(_01919_),
    .X(_01996_));
 sky130_fd_sc_hd__nor2_1 _17707_ (.A(_08404_),
    .B(_09363_),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_1 _17708_ (.A(_10315_),
    .B(_09243_),
    .Y(_01998_));
 sky130_fd_sc_hd__xnor2_1 _17709_ (.A(_01997_),
    .B(_01998_),
    .Y(_01999_));
 sky130_fd_sc_hd__nor2_1 _17710_ (.A(_09647_),
    .B(_09621_),
    .Y(_02000_));
 sky130_fd_sc_hd__xor2_1 _17711_ (.A(_01999_),
    .B(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__o31a_1 _17712_ (.A1(_10059_),
    .A2(_09243_),
    .A3(_01776_),
    .B1(_01887_),
    .X(_02002_));
 sky130_fd_sc_hd__xor2_1 _17713_ (.A(_02001_),
    .B(_02002_),
    .X(_02003_));
 sky130_fd_sc_hd__and2_1 _17714_ (.A(_09519_),
    .B(_09890_),
    .X(_02004_));
 sky130_fd_sc_hd__xor2_1 _17715_ (.A(_02003_),
    .B(_02004_),
    .X(_02005_));
 sky130_fd_sc_hd__o21ai_1 _17716_ (.A1(_01897_),
    .A2(_01903_),
    .B1(_01902_),
    .Y(_02006_));
 sky130_fd_sc_hd__nand2_1 _17717_ (.A(\rbzero.wall_tracer.visualWallDist[4] ),
    .B(_08421_),
    .Y(_02007_));
 sky130_fd_sc_hd__or3_1 _17718_ (.A(_09662_),
    .B(_02007_),
    .C(_01901_),
    .X(_02008_));
 sky130_fd_sc_hd__nor2_1 _17719_ (.A(_09662_),
    .B(_02007_),
    .Y(_02009_));
 sky130_fd_sc_hd__a21o_1 _17720_ (.A1(\rbzero.wall_tracer.visualWallDist[5] ),
    .A2(_01699_),
    .B1(_02009_),
    .X(_02010_));
 sky130_fd_sc_hd__nand2_1 _17721_ (.A(_02008_),
    .B(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__nand2_2 _17722_ (.A(\rbzero.wall_tracer.visualWallDist[6] ),
    .B(_08421_),
    .Y(_02012_));
 sky130_fd_sc_hd__nor2_1 _17723_ (.A(_08428_),
    .B(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__xor2_1 _17724_ (.A(_02011_),
    .B(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__a21bo_1 _17725_ (.A1(_01809_),
    .A2(_01923_),
    .B1_N(_01925_),
    .X(_02015_));
 sky130_fd_sc_hd__and2b_1 _17726_ (.A_N(_02014_),
    .B(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__and2b_1 _17727_ (.A_N(_02015_),
    .B(_02014_),
    .X(_02017_));
 sky130_fd_sc_hd__nor2_1 _17728_ (.A(_02016_),
    .B(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__xnor2_1 _17729_ (.A(_02006_),
    .B(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__a21oi_1 _17730_ (.A1(_01894_),
    .A2(_01907_),
    .B1(_01905_),
    .Y(_02020_));
 sky130_fd_sc_hd__nor2_1 _17731_ (.A(_02019_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__and2_1 _17732_ (.A(_02019_),
    .B(_02020_),
    .X(_02022_));
 sky130_fd_sc_hd__nor2_1 _17733_ (.A(_02021_),
    .B(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__xnor2_1 _17734_ (.A(_02005_),
    .B(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__a21o_1 _17735_ (.A1(_01937_),
    .A2(_01996_),
    .B1(_02024_),
    .X(_02025_));
 sky130_fd_sc_hd__nand3_1 _17736_ (.A(_01937_),
    .B(_01996_),
    .C(_02024_),
    .Y(_02026_));
 sky130_fd_sc_hd__nand2_1 _17737_ (.A(_02025_),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__xnor2_1 _17738_ (.A(_01995_),
    .B(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__or2_1 _17739_ (.A(_09542_),
    .B(_01943_),
    .X(_02029_));
 sky130_fd_sc_hd__or2_1 _17740_ (.A(_01718_),
    .B(_02029_),
    .X(_02030_));
 sky130_fd_sc_hd__nor2_1 _17741_ (.A(_09542_),
    .B(_10093_),
    .Y(_02031_));
 sky130_fd_sc_hd__mux2_1 _17742_ (.A0(_09542_),
    .A1(_02031_),
    .S(_01943_),
    .X(_02032_));
 sky130_fd_sc_hd__xnor2_2 _17743_ (.A(_01831_),
    .B(_02032_),
    .Y(_02033_));
 sky130_fd_sc_hd__a21o_1 _17744_ (.A1(_01832_),
    .A2(_02030_),
    .B1(_02033_),
    .X(_02034_));
 sky130_fd_sc_hd__nand3_1 _17745_ (.A(_01832_),
    .B(_02030_),
    .C(_02033_),
    .Y(_02035_));
 sky130_fd_sc_hd__and2_1 _17746_ (.A(_02034_),
    .B(_02035_),
    .X(_02036_));
 sky130_fd_sc_hd__xnor2_1 _17747_ (.A(_01842_),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__a21boi_1 _17748_ (.A1(_01842_),
    .A2(_01949_),
    .B1_N(_01839_),
    .Y(_02038_));
 sky130_fd_sc_hd__nor2_1 _17749_ (.A(_02037_),
    .B(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__and2_1 _17750_ (.A(_02037_),
    .B(_02038_),
    .X(_02040_));
 sky130_fd_sc_hd__nor2_1 _17751_ (.A(_02039_),
    .B(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__a21o_1 _17752_ (.A1(_01927_),
    .A2(_01935_),
    .B1(_01933_),
    .X(_02042_));
 sky130_fd_sc_hd__a21o_1 _17753_ (.A1(_01941_),
    .A2(_01948_),
    .B1(_01946_),
    .X(_02043_));
 sky130_fd_sc_hd__nor2_1 _17754_ (.A(_10288_),
    .B(_09195_),
    .Y(_02044_));
 sky130_fd_sc_hd__o22a_1 _17755_ (.A1(_10288_),
    .A2(_09315_),
    .B1(_09195_),
    .B2(_01697_),
    .X(_02045_));
 sky130_fd_sc_hd__a21o_1 _17756_ (.A1(_01923_),
    .A2(_02044_),
    .B1(_02045_),
    .X(_02046_));
 sky130_fd_sc_hd__or3_1 _17757_ (.A(_09670_),
    .B(_01922_),
    .C(_02046_),
    .X(_02047_));
 sky130_fd_sc_hd__o21ai_1 _17758_ (.A1(_09670_),
    .A2(_01922_),
    .B1(_02046_),
    .Y(_02048_));
 sky130_fd_sc_hd__and2_1 _17759_ (.A(_02047_),
    .B(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__or2_1 _17760_ (.A(_09528_),
    .B(_01718_),
    .X(_02050_));
 sky130_fd_sc_hd__o22a_1 _17761_ (.A1(_09528_),
    .A2(_10215_),
    .B1(_01718_),
    .B2(_08814_),
    .X(_02051_));
 sky130_fd_sc_hd__o21ba_1 _17762_ (.A1(_01928_),
    .A2(_02050_),
    .B1_N(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__nor2_1 _17763_ (.A(_01818_),
    .B(_09560_),
    .Y(_02053_));
 sky130_fd_sc_hd__xnor2_1 _17764_ (.A(_02052_),
    .B(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__or3_1 _17765_ (.A(_01818_),
    .B(_09677_),
    .C(_01929_),
    .X(_02055_));
 sky130_fd_sc_hd__o21a_1 _17766_ (.A1(_01814_),
    .A2(_01928_),
    .B1(_02055_),
    .X(_02056_));
 sky130_fd_sc_hd__xor2_1 _17767_ (.A(_02054_),
    .B(_02056_),
    .X(_02057_));
 sky130_fd_sc_hd__xnor2_1 _17768_ (.A(_02049_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__xor2_1 _17769_ (.A(_02043_),
    .B(_02058_),
    .X(_02059_));
 sky130_fd_sc_hd__xnor2_1 _17770_ (.A(_02042_),
    .B(_02059_),
    .Y(_02060_));
 sky130_fd_sc_hd__xnor2_1 _17771_ (.A(_02041_),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__a21oi_1 _17772_ (.A1(_01940_),
    .A2(_01954_),
    .B1(_01952_),
    .Y(_02062_));
 sky130_fd_sc_hd__nor2_1 _17773_ (.A(_02061_),
    .B(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__and2_1 _17774_ (.A(_02061_),
    .B(_02062_),
    .X(_02064_));
 sky130_fd_sc_hd__nor2_1 _17775_ (.A(_02063_),
    .B(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__xnor2_1 _17776_ (.A(_02028_),
    .B(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__nor2_1 _17777_ (.A(_01955_),
    .B(_01956_),
    .Y(_02067_));
 sky130_fd_sc_hd__a21oi_1 _17778_ (.A1(_01918_),
    .A2(_01957_),
    .B1(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__xor2_1 _17779_ (.A(_02066_),
    .B(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__xnor2_1 _17780_ (.A(_01994_),
    .B(_02069_),
    .Y(_02070_));
 sky130_fd_sc_hd__nor2_1 _17781_ (.A(_01958_),
    .B(_01960_),
    .Y(_02071_));
 sky130_fd_sc_hd__a21oi_1 _17782_ (.A1(_01880_),
    .A2(_01961_),
    .B1(_02071_),
    .Y(_02072_));
 sky130_fd_sc_hd__nor2_1 _17783_ (.A(_02070_),
    .B(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__and2_1 _17784_ (.A(_02070_),
    .B(_02072_),
    .X(_02074_));
 sky130_fd_sc_hd__nor2_1 _17785_ (.A(_02073_),
    .B(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__xnor2_1 _17786_ (.A(_01878_),
    .B(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__a21o_1 _17787_ (.A1(_01965_),
    .A2(_01968_),
    .B1(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__and3_2 _17788_ (.A(_01965_),
    .B(_01968_),
    .C(_02076_),
    .X(_02078_));
 sky130_fd_sc_hd__inv_2 _17789_ (.A(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__nand2_1 _17790_ (.A(_02077_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__a21oi_1 _17791_ (.A1(_01972_),
    .A2(_01980_),
    .B1(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__a31o_1 _17792_ (.A1(_01972_),
    .A2(_01980_),
    .A3(_02080_),
    .B1(_08123_),
    .X(_02082_));
 sky130_fd_sc_hd__or2_1 _17793_ (.A(_02081_),
    .B(_02082_),
    .X(_02083_));
 sky130_fd_sc_hd__o21ai_1 _17794_ (.A1(_01988_),
    .A2(_01989_),
    .B1(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__mux2_1 _17795_ (.A0(\rbzero.wall_tracer.trackDistX[7] ),
    .A1(_02084_),
    .S(_09844_),
    .X(_02085_));
 sky130_fd_sc_hd__clkbuf_1 _17796_ (.A(_02085_),
    .X(_00546_));
 sky130_fd_sc_hd__or2b_1 _17797_ (.A(_02027_),
    .B_N(_01995_),
    .X(_02086_));
 sky130_fd_sc_hd__o2bb2a_1 _17798_ (.A1_N(_02003_),
    .A2_N(_02004_),
    .B1(_02001_),
    .B2(_02002_),
    .X(_02087_));
 sky130_fd_sc_hd__a21o_1 _17799_ (.A1(_02025_),
    .A2(_02086_),
    .B1(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__nand3_1 _17800_ (.A(_02025_),
    .B(_02086_),
    .C(_02087_),
    .Y(_02089_));
 sky130_fd_sc_hd__and2_1 _17801_ (.A(_02088_),
    .B(_02089_),
    .X(_02090_));
 sky130_fd_sc_hd__a21bo_1 _17802_ (.A1(_01842_),
    .A2(_02036_),
    .B1_N(_01839_),
    .X(_02091_));
 sky130_fd_sc_hd__and2_1 _17803_ (.A(_01832_),
    .B(_02029_),
    .X(_02092_));
 sky130_fd_sc_hd__xor2_2 _17804_ (.A(_02033_),
    .B(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__xor2_1 _17805_ (.A(_01842_),
    .B(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__xor2_1 _17806_ (.A(_02091_),
    .B(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__nand2_1 _17807_ (.A(_02049_),
    .B(_02057_),
    .Y(_02096_));
 sky130_fd_sc_hd__o21ai_1 _17808_ (.A1(_02054_),
    .A2(_02056_),
    .B1(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__nand2_1 _17809_ (.A(_01831_),
    .B(_02032_),
    .Y(_02098_));
 sky130_fd_sc_hd__nand2_1 _17810_ (.A(_02098_),
    .B(_02034_),
    .Y(_02099_));
 sky130_fd_sc_hd__nor2_1 _17811_ (.A(_01697_),
    .B(_09433_),
    .Y(_02100_));
 sky130_fd_sc_hd__xnor2_1 _17812_ (.A(_02044_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__or3_1 _17813_ (.A(_01922_),
    .B(_09315_),
    .C(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__o21ai_1 _17814_ (.A1(_01922_),
    .A2(_09315_),
    .B1(_02101_),
    .Y(_02103_));
 sky130_fd_sc_hd__and2_1 _17815_ (.A(_02102_),
    .B(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__nor2_1 _17816_ (.A(_08814_),
    .B(_10093_),
    .Y(_02105_));
 sky130_fd_sc_hd__xnor2_1 _17817_ (.A(_02050_),
    .B(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__nor2_1 _17818_ (.A(_01818_),
    .B(_10215_),
    .Y(_02107_));
 sky130_fd_sc_hd__xnor2_1 _17819_ (.A(_02106_),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__o32a_1 _17820_ (.A1(_01818_),
    .A2(_09560_),
    .A3(_02051_),
    .B1(_02050_),
    .B2(_01928_),
    .X(_02109_));
 sky130_fd_sc_hd__nor2_1 _17821_ (.A(_02108_),
    .B(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__and2_1 _17822_ (.A(_02108_),
    .B(_02109_),
    .X(_02111_));
 sky130_fd_sc_hd__nor2_1 _17823_ (.A(_02110_),
    .B(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__xor2_1 _17824_ (.A(_02104_),
    .B(_02112_),
    .X(_02113_));
 sky130_fd_sc_hd__xnor2_1 _17825_ (.A(_02099_),
    .B(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__xnor2_1 _17826_ (.A(_02097_),
    .B(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__and2_1 _17827_ (.A(_02095_),
    .B(_02115_),
    .X(_02116_));
 sky130_fd_sc_hd__nor2_1 _17828_ (.A(_02095_),
    .B(_02115_),
    .Y(_02117_));
 sky130_fd_sc_hd__or2_1 _17829_ (.A(_02116_),
    .B(_02117_),
    .X(_02118_));
 sky130_fd_sc_hd__a21oi_1 _17830_ (.A1(_02041_),
    .A2(_02060_),
    .B1(_02039_),
    .Y(_02119_));
 sky130_fd_sc_hd__xor2_1 _17831_ (.A(_02118_),
    .B(_02119_),
    .X(_02120_));
 sky130_fd_sc_hd__a21o_1 _17832_ (.A1(_02005_),
    .A2(_02023_),
    .B1(_02021_),
    .X(_02121_));
 sky130_fd_sc_hd__or2b_1 _17833_ (.A(_02058_),
    .B_N(_02043_),
    .X(_02122_));
 sky130_fd_sc_hd__or2b_1 _17834_ (.A(_02059_),
    .B_N(_02042_),
    .X(_02123_));
 sky130_fd_sc_hd__or2_1 _17835_ (.A(_08499_),
    .B(_09243_),
    .X(_02124_));
 sky130_fd_sc_hd__or3_1 _17836_ (.A(_10315_),
    .B(_09363_),
    .C(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__o21ai_1 _17837_ (.A1(_10315_),
    .A2(_09363_),
    .B1(_02124_),
    .Y(_02126_));
 sky130_fd_sc_hd__nand2_1 _17838_ (.A(_02125_),
    .B(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__nor2_1 _17839_ (.A(_10059_),
    .B(_09621_),
    .Y(_02128_));
 sky130_fd_sc_hd__xor2_1 _17840_ (.A(_02127_),
    .B(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__nand2_1 _17841_ (.A(_01997_),
    .B(_01998_),
    .Y(_02130_));
 sky130_fd_sc_hd__o31a_1 _17842_ (.A1(_09647_),
    .A2(_09621_),
    .A3(_01999_),
    .B1(_02130_),
    .X(_02131_));
 sky130_fd_sc_hd__xor2_1 _17843_ (.A(_02129_),
    .B(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__and2_1 _17844_ (.A(_09647_),
    .B(_09890_),
    .X(_02133_));
 sky130_fd_sc_hd__xor2_1 _17845_ (.A(_02132_),
    .B(_02133_),
    .X(_02134_));
 sky130_fd_sc_hd__o31ai_2 _17846_ (.A1(_08428_),
    .A2(_02012_),
    .A3(_02011_),
    .B1(_02008_),
    .Y(_02135_));
 sky130_fd_sc_hd__nand2_1 _17847_ (.A(_01923_),
    .B(_02044_),
    .Y(_02136_));
 sky130_fd_sc_hd__nor2_1 _17848_ (.A(_09670_),
    .B(_01898_),
    .Y(_02137_));
 sky130_fd_sc_hd__nand2_1 _17849_ (.A(_02009_),
    .B(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__o22ai_1 _17850_ (.A1(_09670_),
    .A2(_02007_),
    .B1(_01898_),
    .B2(_09662_),
    .Y(_02139_));
 sky130_fd_sc_hd__nand2_1 _17851_ (.A(_02138_),
    .B(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__nor2_1 _17852_ (.A(_08476_),
    .B(_02012_),
    .Y(_02141_));
 sky130_fd_sc_hd__xor2_1 _17853_ (.A(_02140_),
    .B(_02141_),
    .X(_02142_));
 sky130_fd_sc_hd__a21oi_1 _17854_ (.A1(_02136_),
    .A2(_02047_),
    .B1(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__and3_1 _17855_ (.A(_02136_),
    .B(_02047_),
    .C(_02142_),
    .X(_02144_));
 sky130_fd_sc_hd__nor2_1 _17856_ (.A(_02143_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__xnor2_1 _17857_ (.A(_02135_),
    .B(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hd__a21oi_1 _17858_ (.A1(_02006_),
    .A2(_02018_),
    .B1(_02016_),
    .Y(_02147_));
 sky130_fd_sc_hd__nor2_1 _17859_ (.A(_02146_),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__and2_1 _17860_ (.A(_02146_),
    .B(_02147_),
    .X(_02149_));
 sky130_fd_sc_hd__nor2_1 _17861_ (.A(_02148_),
    .B(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__xnor2_1 _17862_ (.A(_02134_),
    .B(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__a21o_1 _17863_ (.A1(_02122_),
    .A2(_02123_),
    .B1(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__nand3_1 _17864_ (.A(_02122_),
    .B(_02123_),
    .C(_02151_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2_1 _17865_ (.A(_02152_),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__xnor2_1 _17866_ (.A(_02121_),
    .B(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_1 _17867_ (.A(_02120_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__or2_1 _17868_ (.A(_02120_),
    .B(_02155_),
    .X(_02157_));
 sky130_fd_sc_hd__nand2_1 _17869_ (.A(_02156_),
    .B(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__a21oi_1 _17870_ (.A1(_02028_),
    .A2(_02065_),
    .B1(_02063_),
    .Y(_02159_));
 sky130_fd_sc_hd__xor2_1 _17871_ (.A(_02158_),
    .B(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__nand2_1 _17872_ (.A(_02090_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__or2_1 _17873_ (.A(_02090_),
    .B(_02160_),
    .X(_02162_));
 sky130_fd_sc_hd__nand2_1 _17874_ (.A(_02161_),
    .B(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__nor2_1 _17875_ (.A(_02066_),
    .B(_02068_),
    .Y(_02164_));
 sky130_fd_sc_hd__a21oi_2 _17876_ (.A1(_01994_),
    .A2(_02069_),
    .B1(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__xor2_1 _17877_ (.A(_02163_),
    .B(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__xnor2_1 _17878_ (.A(_01992_),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__a21oi_2 _17879_ (.A1(_01878_),
    .A2(_02075_),
    .B1(_02073_),
    .Y(_02168_));
 sky130_fd_sc_hd__or2_1 _17880_ (.A(_02167_),
    .B(_02168_),
    .X(_02169_));
 sky130_fd_sc_hd__nand2_1 _17881_ (.A(_02167_),
    .B(_02168_),
    .Y(_02170_));
 sky130_fd_sc_hd__and2_1 _17882_ (.A(_02169_),
    .B(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__inv_2 _17883_ (.A(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__a311o_1 _17884_ (.A1(_01972_),
    .A2(_01980_),
    .A3(_02077_),
    .B1(_02078_),
    .C1(_02172_),
    .X(_02173_));
 sky130_fd_sc_hd__a31o_1 _17885_ (.A1(_01972_),
    .A2(_01980_),
    .A3(_02077_),
    .B1(_02078_),
    .X(_02174_));
 sky130_fd_sc_hd__a21oi_1 _17886_ (.A1(_02172_),
    .A2(_02174_),
    .B1(_08124_),
    .Y(_02175_));
 sky130_fd_sc_hd__nand2_1 _17887_ (.A(_02173_),
    .B(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__or2_1 _17888_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .X(_02177_));
 sky130_fd_sc_hd__nand2_1 _17889_ (.A(\rbzero.wall_tracer.trackDistX[8] ),
    .B(\rbzero.wall_tracer.stepDistX[8] ),
    .Y(_02178_));
 sky130_fd_sc_hd__nand2_1 _17890_ (.A(_02177_),
    .B(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__o21a_1 _17891_ (.A1(_01984_),
    .A2(_01987_),
    .B1(_01985_),
    .X(_02180_));
 sky130_fd_sc_hd__or2_1 _17892_ (.A(_02179_),
    .B(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__a21oi_1 _17893_ (.A1(_02179_),
    .A2(_02180_),
    .B1(_06105_),
    .Y(_02182_));
 sky130_fd_sc_hd__a21oi_1 _17894_ (.A1(_02181_),
    .A2(_02182_),
    .B1(_09785_),
    .Y(_02183_));
 sky130_fd_sc_hd__o2bb2a_1 _17895_ (.A1_N(_02176_),
    .A2_N(_02183_),
    .B1(\rbzero.wall_tracer.trackDistX[8] ),
    .B2(_09879_),
    .X(_00547_));
 sky130_fd_sc_hd__or2_1 _17896_ (.A(_02163_),
    .B(_02165_),
    .X(_02184_));
 sky130_fd_sc_hd__nand2_1 _17897_ (.A(_01992_),
    .B(_02166_),
    .Y(_02185_));
 sky130_fd_sc_hd__and2_1 _17898_ (.A(_02091_),
    .B(_02094_),
    .X(_02186_));
 sky130_fd_sc_hd__a21o_1 _17899_ (.A1(_02104_),
    .A2(_02112_),
    .B1(_02110_),
    .X(_02187_));
 sky130_fd_sc_hd__o21a_1 _17900_ (.A1(_02033_),
    .A2(_02092_),
    .B1(_02098_),
    .X(_02188_));
 sky130_fd_sc_hd__nor2_1 _17901_ (.A(_01697_),
    .B(_10214_),
    .Y(_02189_));
 sky130_fd_sc_hd__nor2_1 _17902_ (.A(_10288_),
    .B(_09433_),
    .Y(_02190_));
 sky130_fd_sc_hd__xnor2_1 _17903_ (.A(_02189_),
    .B(_02190_),
    .Y(_02191_));
 sky130_fd_sc_hd__or2_1 _17904_ (.A(_01922_),
    .B(_09195_),
    .X(_02192_));
 sky130_fd_sc_hd__xnor2_1 _17905_ (.A(_02191_),
    .B(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__nand2_1 _17906_ (.A(_08530_),
    .B(_02105_),
    .Y(_02194_));
 sky130_fd_sc_hd__a2bb2o_1 _17907_ (.A1_N(_01718_),
    .A2_N(_02194_),
    .B1(_02106_),
    .B2(_02107_),
    .X(_02195_));
 sky130_fd_sc_hd__a21o_1 _17908_ (.A1(_08814_),
    .A2(_09528_),
    .B1(_10093_),
    .X(_02196_));
 sky130_fd_sc_hd__a21o_1 _17909_ (.A1(_08530_),
    .A2(_02105_),
    .B1(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__nor2_1 _17910_ (.A(_01818_),
    .B(_01718_),
    .Y(_02198_));
 sky130_fd_sc_hd__xnor2_1 _17911_ (.A(_02197_),
    .B(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__xor2_1 _17912_ (.A(_02195_),
    .B(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__xnor2_1 _17913_ (.A(_02193_),
    .B(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__and2b_1 _17914_ (.A_N(_02188_),
    .B(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__and2b_1 _17915_ (.A_N(_02201_),
    .B(_02188_),
    .X(_02203_));
 sky130_fd_sc_hd__nor2_1 _17916_ (.A(_02202_),
    .B(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__xnor2_1 _17917_ (.A(_02187_),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__and3_1 _17918_ (.A(_10221_),
    .B(_01729_),
    .C(_02093_),
    .X(_02206_));
 sky130_fd_sc_hd__o22a_1 _17919_ (.A1(_01840_),
    .A2(_02093_),
    .B1(_02205_),
    .B2(_02206_),
    .X(_02207_));
 sky130_fd_sc_hd__nor3_1 _17920_ (.A(_01840_),
    .B(_02093_),
    .C(_02205_),
    .Y(_02208_));
 sky130_fd_sc_hd__o2bb2a_1 _17921_ (.A1_N(_02205_),
    .A2_N(_02206_),
    .B1(_02207_),
    .B2(_02208_),
    .X(_02209_));
 sky130_fd_sc_hd__o21a_1 _17922_ (.A1(_02186_),
    .A2(_02116_),
    .B1(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__nor3_1 _17923_ (.A(_02186_),
    .B(_02116_),
    .C(_02209_),
    .Y(_02211_));
 sky130_fd_sc_hd__nor2_1 _17924_ (.A(_02210_),
    .B(_02211_),
    .Y(_02212_));
 sky130_fd_sc_hd__a21o_1 _17925_ (.A1(_02134_),
    .A2(_02150_),
    .B1(_02148_),
    .X(_02213_));
 sky130_fd_sc_hd__or2b_1 _17926_ (.A(_02114_),
    .B_N(_02097_),
    .X(_02214_));
 sky130_fd_sc_hd__a21bo_1 _17927_ (.A1(_02099_),
    .A2(_02113_),
    .B1_N(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__nand2_1 _17928_ (.A(\rbzero.wall_tracer.visualWallDist[8] ),
    .B(_01699_),
    .Y(_02216_));
 sky130_fd_sc_hd__a22o_1 _17929_ (.A1(\rbzero.wall_tracer.visualWallDist[8] ),
    .A2(_10183_),
    .B1(_01699_),
    .B2(\rbzero.wall_tracer.visualWallDist[7] ),
    .X(_02217_));
 sky130_fd_sc_hd__o21ai_1 _17930_ (.A1(_02124_),
    .A2(_02216_),
    .B1(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__or3_1 _17931_ (.A(_10315_),
    .B(_09621_),
    .C(_02218_),
    .X(_02219_));
 sky130_fd_sc_hd__o21ai_1 _17932_ (.A1(_10315_),
    .A2(_09621_),
    .B1(_02218_),
    .Y(_02220_));
 sky130_fd_sc_hd__nand2_1 _17933_ (.A(_02219_),
    .B(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__o31a_1 _17934_ (.A1(_10059_),
    .A2(_09621_),
    .A3(_02127_),
    .B1(_02125_),
    .X(_02222_));
 sky130_fd_sc_hd__xnor2_1 _17935_ (.A(_02221_),
    .B(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__nand2_1 _17936_ (.A(_10059_),
    .B(_09890_),
    .Y(_02224_));
 sky130_fd_sc_hd__xnor2_1 _17937_ (.A(_02223_),
    .B(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__a21bo_1 _17938_ (.A1(_02139_),
    .A2(_02141_),
    .B1_N(_02138_),
    .X(_02226_));
 sky130_fd_sc_hd__a21bo_1 _17939_ (.A1(_02044_),
    .A2(_02100_),
    .B1_N(_02102_),
    .X(_02227_));
 sky130_fd_sc_hd__nor2_1 _17940_ (.A(_02007_),
    .B(_09315_),
    .Y(_02228_));
 sky130_fd_sc_hd__xnor2_1 _17941_ (.A(_02137_),
    .B(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__nor2_1 _17942_ (.A(_09662_),
    .B(_02012_),
    .Y(_02230_));
 sky130_fd_sc_hd__xnor2_1 _17943_ (.A(_02229_),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__xor2_1 _17944_ (.A(_02227_),
    .B(_02231_),
    .X(_02232_));
 sky130_fd_sc_hd__and2_1 _17945_ (.A(_02226_),
    .B(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__nor2_1 _17946_ (.A(_02226_),
    .B(_02232_),
    .Y(_02234_));
 sky130_fd_sc_hd__or2_1 _17947_ (.A(_02233_),
    .B(_02234_),
    .X(_02235_));
 sky130_fd_sc_hd__a21oi_1 _17948_ (.A1(_02135_),
    .A2(_02145_),
    .B1(_02143_),
    .Y(_02236_));
 sky130_fd_sc_hd__or2_1 _17949_ (.A(_02235_),
    .B(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__nand2_1 _17950_ (.A(_02235_),
    .B(_02236_),
    .Y(_02238_));
 sky130_fd_sc_hd__and2_1 _17951_ (.A(_02237_),
    .B(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__xnor2_1 _17952_ (.A(_02225_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__xnor2_1 _17953_ (.A(_02215_),
    .B(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__xnor2_1 _17954_ (.A(_02213_),
    .B(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__xnor2_1 _17955_ (.A(_02212_),
    .B(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__o21a_1 _17956_ (.A1(_02118_),
    .A2(_02119_),
    .B1(_02156_),
    .X(_02244_));
 sky130_fd_sc_hd__xnor2_1 _17957_ (.A(_02243_),
    .B(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__or2b_1 _17958_ (.A(_02154_),
    .B_N(_02121_),
    .X(_02246_));
 sky130_fd_sc_hd__o2bb2a_1 _17959_ (.A1_N(_02132_),
    .A2_N(_02133_),
    .B1(_02129_),
    .B2(_02131_),
    .X(_02247_));
 sky130_fd_sc_hd__a21o_1 _17960_ (.A1(_02152_),
    .A2(_02246_),
    .B1(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__nand3_1 _17961_ (.A(_02152_),
    .B(_02246_),
    .C(_02247_),
    .Y(_02249_));
 sky130_fd_sc_hd__and2_1 _17962_ (.A(_02248_),
    .B(_02249_),
    .X(_02250_));
 sky130_fd_sc_hd__xor2_1 _17963_ (.A(_02245_),
    .B(_02250_),
    .X(_02251_));
 sky130_fd_sc_hd__o21a_1 _17964_ (.A1(_02158_),
    .A2(_02159_),
    .B1(_02161_),
    .X(_02252_));
 sky130_fd_sc_hd__xor2_1 _17965_ (.A(_02251_),
    .B(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__xor2_1 _17966_ (.A(_02088_),
    .B(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__a21o_1 _17967_ (.A1(_02184_),
    .A2(_02185_),
    .B1(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__inv_2 _17968_ (.A(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__and3_1 _17969_ (.A(_02184_),
    .B(_02185_),
    .C(_02254_),
    .X(_02257_));
 sky130_fd_sc_hd__nor2_1 _17970_ (.A(_02256_),
    .B(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__inv_2 _17971_ (.A(_02258_),
    .Y(_02259_));
 sky130_fd_sc_hd__a21oi_1 _17972_ (.A1(_02169_),
    .A2(_02173_),
    .B1(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__a31o_1 _17973_ (.A1(_02169_),
    .A2(_02173_),
    .A3(_02259_),
    .B1(_01757_),
    .X(_02261_));
 sky130_fd_sc_hd__or2_1 _17974_ (.A(_02260_),
    .B(_02261_),
    .X(_02262_));
 sky130_fd_sc_hd__and2_1 _17975_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .X(_02263_));
 sky130_fd_sc_hd__nor2_1 _17976_ (.A(\rbzero.wall_tracer.trackDistX[9] ),
    .B(\rbzero.wall_tracer.stepDistX[9] ),
    .Y(_02264_));
 sky130_fd_sc_hd__nor2_1 _17977_ (.A(_02263_),
    .B(_02264_),
    .Y(_02265_));
 sky130_fd_sc_hd__nand2_1 _17978_ (.A(_02178_),
    .B(_02180_),
    .Y(_02266_));
 sky130_fd_sc_hd__and2_1 _17979_ (.A(_02177_),
    .B(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__xnor2_1 _17980_ (.A(_02265_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__o21a_1 _17981_ (.A1(_09872_),
    .A2(_02268_),
    .B1(_09879_),
    .X(_02269_));
 sky130_fd_sc_hd__o2bb2a_1 _17982_ (.A1_N(_02262_),
    .A2_N(_02269_),
    .B1(\rbzero.wall_tracer.trackDistX[9] ),
    .B2(_09879_),
    .X(_00548_));
 sky130_fd_sc_hd__a21o_1 _17983_ (.A1(_02169_),
    .A2(_02255_),
    .B1(_02257_),
    .X(_02270_));
 sky130_fd_sc_hd__or2b_1 _17984_ (.A(_02088_),
    .B_N(_02253_),
    .X(_02271_));
 sky130_fd_sc_hd__o21ai_1 _17985_ (.A1(_02251_),
    .A2(_02252_),
    .B1(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__o22a_1 _17986_ (.A1(_02221_),
    .A2(_02222_),
    .B1(_02223_),
    .B2(_02224_),
    .X(_02273_));
 sky130_fd_sc_hd__o21a_1 _17987_ (.A1(_02196_),
    .A2(_02198_),
    .B1(_02194_),
    .X(_02274_));
 sky130_fd_sc_hd__and2b_1 _17988_ (.A_N(_02241_),
    .B(_02213_),
    .X(_02275_));
 sky130_fd_sc_hd__a21oi_1 _17989_ (.A1(_02215_),
    .A2(_02240_),
    .B1(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__xnor2_1 _17990_ (.A(_02274_),
    .B(_02276_),
    .Y(_02277_));
 sky130_fd_sc_hd__xor2_1 _17991_ (.A(_02188_),
    .B(_02207_),
    .X(_02278_));
 sky130_fd_sc_hd__a21oi_1 _17992_ (.A1(_02187_),
    .A2(_02204_),
    .B1(_02202_),
    .Y(_02279_));
 sky130_fd_sc_hd__nand2_1 _17993_ (.A(_02189_),
    .B(_02190_),
    .Y(_02280_));
 sky130_fd_sc_hd__o31a_1 _17994_ (.A1(_01922_),
    .A2(_09195_),
    .A3(_02191_),
    .B1(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__o21a_1 _17995_ (.A1(_02124_),
    .A2(_02216_),
    .B1(_02219_),
    .X(_02282_));
 sky130_fd_sc_hd__nor2_1 _17996_ (.A(_08499_),
    .B(_09621_),
    .Y(_02283_));
 sky130_fd_sc_hd__xnor2_1 _17997_ (.A(_02282_),
    .B(_02283_),
    .Y(_02284_));
 sky130_fd_sc_hd__xnor2_1 _17998_ (.A(_02281_),
    .B(_02284_),
    .Y(_02285_));
 sky130_fd_sc_hd__nand2_1 _17999_ (.A(_02137_),
    .B(_02228_),
    .Y(_02286_));
 sky130_fd_sc_hd__o31a_1 _18000_ (.A1(_09662_),
    .A2(_02012_),
    .A3(_02229_),
    .B1(_02286_),
    .X(_02287_));
 sky130_fd_sc_hd__nor2_1 _18001_ (.A(_09670_),
    .B(_02012_),
    .Y(_02288_));
 sky130_fd_sc_hd__xnor2_1 _18002_ (.A(_02287_),
    .B(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__nor2_1 _18003_ (.A(_08455_),
    .B(_09243_),
    .Y(_02290_));
 sky130_fd_sc_hd__xnor2_1 _18004_ (.A(_02216_),
    .B(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__xnor2_1 _18005_ (.A(_02289_),
    .B(_02291_),
    .Y(_02292_));
 sky130_fd_sc_hd__xnor2_1 _18006_ (.A(_02285_),
    .B(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__xnor2_1 _18007_ (.A(_02279_),
    .B(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__xnor2_1 _18008_ (.A(_02278_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__xnor2_1 _18009_ (.A(_02277_),
    .B(_02295_),
    .Y(_02296_));
 sky130_fd_sc_hd__a21o_1 _18010_ (.A1(_02212_),
    .A2(_02242_),
    .B1(_02210_),
    .X(_02297_));
 sky130_fd_sc_hd__and2b_1 _18011_ (.A_N(_02193_),
    .B(_02200_),
    .X(_02298_));
 sky130_fd_sc_hd__a21o_1 _18012_ (.A1(_02195_),
    .A2(_02199_),
    .B1(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__nor2_1 _18013_ (.A(_01922_),
    .B(_09433_),
    .Y(_02300_));
 sky130_fd_sc_hd__xnor2_1 _18014_ (.A(_02299_),
    .B(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__or2b_1 _18015_ (.A(_02225_),
    .B_N(_02239_),
    .X(_02302_));
 sky130_fd_sc_hd__a21oi_1 _18016_ (.A1(_02227_),
    .A2(_02231_),
    .B1(_02233_),
    .Y(_02303_));
 sky130_fd_sc_hd__o211a_1 _18017_ (.A1(_09315_),
    .A2(_01898_),
    .B1(_09890_),
    .C1(_10315_),
    .X(_02304_));
 sky130_fd_sc_hd__a211oi_1 _18018_ (.A1(_10315_),
    .A2(_09890_),
    .B1(_01898_),
    .C1(_09315_),
    .Y(_02305_));
 sky130_fd_sc_hd__nor2_1 _18019_ (.A(_02304_),
    .B(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__xnor2_1 _18020_ (.A(_02303_),
    .B(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__a21oi_1 _18021_ (.A1(_02237_),
    .A2(_02302_),
    .B1(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__a31o_1 _18022_ (.A1(_02237_),
    .A2(_02302_),
    .A3(_02307_),
    .B1(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__nor2_1 _18023_ (.A(_01818_),
    .B(_10093_),
    .Y(_02310_));
 sky130_fd_sc_hd__nor2_1 _18024_ (.A(_10288_),
    .B(_10214_),
    .Y(_02311_));
 sky130_fd_sc_hd__nor2_1 _18025_ (.A(_01697_),
    .B(_09974_),
    .Y(_02312_));
 sky130_fd_sc_hd__xor2_1 _18026_ (.A(_02311_),
    .B(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__xnor2_1 _18027_ (.A(_02310_),
    .B(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__nor2_1 _18028_ (.A(_02007_),
    .B(_09195_),
    .Y(_02315_));
 sky130_fd_sc_hd__xnor2_1 _18029_ (.A(_02314_),
    .B(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__xnor2_1 _18030_ (.A(_02309_),
    .B(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__xnor2_1 _18031_ (.A(_02301_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__xnor2_1 _18032_ (.A(_02248_),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__xnor2_1 _18033_ (.A(_02297_),
    .B(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hd__xnor2_1 _18034_ (.A(_02296_),
    .B(_02320_),
    .Y(_02321_));
 sky130_fd_sc_hd__or2b_1 _18035_ (.A(_02245_),
    .B_N(_02250_),
    .X(_02322_));
 sky130_fd_sc_hd__o21a_1 _18036_ (.A1(_02243_),
    .A2(_02244_),
    .B1(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__xnor2_1 _18037_ (.A(_02321_),
    .B(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__xnor2_1 _18038_ (.A(_02273_),
    .B(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__xnor2_1 _18039_ (.A(_02272_),
    .B(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__o211a_1 _18040_ (.A1(_02173_),
    .A2(_02259_),
    .B1(_02270_),
    .C1(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__a311o_1 _18041_ (.A1(_02169_),
    .A2(_02173_),
    .A3(_02255_),
    .B1(_02257_),
    .C1(_02326_),
    .X(_02328_));
 sky130_fd_sc_hd__or3b_1 _18042_ (.A(_08124_),
    .B(_02327_),
    .C_N(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__a31o_1 _18043_ (.A1(_02177_),
    .A2(_02265_),
    .A3(_02266_),
    .B1(_02263_),
    .X(_02330_));
 sky130_fd_sc_hd__xnor2_1 _18044_ (.A(\rbzero.wall_tracer.trackDistX[10] ),
    .B(\rbzero.wall_tracer.stepDistX[10] ),
    .Y(_02331_));
 sky130_fd_sc_hd__xnor2_1 _18045_ (.A(_02330_),
    .B(_02331_),
    .Y(_02332_));
 sky130_fd_sc_hd__a21oi_1 _18046_ (.A1(_08124_),
    .A2(_02332_),
    .B1(_09783_),
    .Y(_02333_));
 sky130_fd_sc_hd__o2bb2a_1 _18047_ (.A1_N(_02329_),
    .A2_N(_02333_),
    .B1(\rbzero.wall_tracer.trackDistX[10] ),
    .B2(_09879_),
    .X(_00549_));
 sky130_fd_sc_hd__and2_1 _18048_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .X(_02334_));
 sky130_fd_sc_hd__nor2_1 _18049_ (.A(\rbzero.wall_tracer.trackDistY[-11] ),
    .B(\rbzero.wall_tracer.stepDistY[-11] ),
    .Y(_02335_));
 sky130_fd_sc_hd__o21a_2 _18050_ (.A1(_08139_),
    .A2(_08405_),
    .B1(_04433_),
    .X(_02336_));
 sky130_fd_sc_hd__buf_4 _18051_ (.A(_02336_),
    .X(_02337_));
 sky130_fd_sc_hd__o31a_1 _18052_ (.A1(_09872_),
    .A2(_02334_),
    .A3(_02335_),
    .B1(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__buf_4 _18053_ (.A(_02336_),
    .X(_02339_));
 sky130_fd_sc_hd__buf_2 _18054_ (.A(_02339_),
    .X(_02340_));
 sky130_fd_sc_hd__o2bb2a_1 _18055_ (.A1_N(_09804_),
    .A2_N(_02338_),
    .B1(_02340_),
    .B2(\rbzero.wall_tracer.trackDistY[-11] ),
    .X(_00550_));
 sky130_fd_sc_hd__clkbuf_4 _18056_ (.A(_06104_),
    .X(_02341_));
 sky130_fd_sc_hd__or2_1 _18057_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .X(_02342_));
 sky130_fd_sc_hd__nand2_1 _18058_ (.A(\rbzero.wall_tracer.trackDistY[-10] ),
    .B(\rbzero.wall_tracer.stepDistY[-10] ),
    .Y(_02343_));
 sky130_fd_sc_hd__and3_1 _18059_ (.A(_02334_),
    .B(_02342_),
    .C(_02343_),
    .X(_02344_));
 sky130_fd_sc_hd__a21oi_1 _18060_ (.A1(_02342_),
    .A2(_02343_),
    .B1(_02334_),
    .Y(_02345_));
 sky130_fd_sc_hd__o31a_1 _18061_ (.A1(_02341_),
    .A2(_02344_),
    .A3(_02345_),
    .B1(_02337_),
    .X(_02346_));
 sky130_fd_sc_hd__o2bb2a_1 _18062_ (.A1_N(_09815_),
    .A2_N(_02346_),
    .B1(_02340_),
    .B2(\rbzero.wall_tracer.trackDistY[-10] ),
    .X(_00551_));
 sky130_fd_sc_hd__a21oi_1 _18063_ (.A1(\rbzero.wall_tracer.trackDistY[-10] ),
    .A2(\rbzero.wall_tracer.stepDistY[-10] ),
    .B1(_02344_),
    .Y(_02347_));
 sky130_fd_sc_hd__nor2_1 _18064_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .Y(_02348_));
 sky130_fd_sc_hd__and2_1 _18065_ (.A(\rbzero.wall_tracer.trackDistY[-9] ),
    .B(\rbzero.wall_tracer.stepDistY[-9] ),
    .X(_02349_));
 sky130_fd_sc_hd__nor3_1 _18066_ (.A(_02347_),
    .B(_02348_),
    .C(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__o21a_1 _18067_ (.A1(_02348_),
    .A2(_02349_),
    .B1(_02347_),
    .X(_02351_));
 sky130_fd_sc_hd__o31a_1 _18068_ (.A1(_02341_),
    .A2(_02350_),
    .A3(_02351_),
    .B1(_02337_),
    .X(_02352_));
 sky130_fd_sc_hd__o2bb2a_1 _18069_ (.A1_N(_09823_),
    .A2_N(_02352_),
    .B1(_02340_),
    .B2(\rbzero.wall_tracer.trackDistY[-9] ),
    .X(_00552_));
 sky130_fd_sc_hd__or2_1 _18070_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .X(_02353_));
 sky130_fd_sc_hd__nand2_1 _18071_ (.A(\rbzero.wall_tracer.trackDistY[-8] ),
    .B(\rbzero.wall_tracer.stepDistY[-8] ),
    .Y(_02354_));
 sky130_fd_sc_hd__o21bai_1 _18072_ (.A1(_02347_),
    .A2(_02348_),
    .B1_N(_02349_),
    .Y(_02355_));
 sky130_fd_sc_hd__and3_1 _18073_ (.A(_02353_),
    .B(_02354_),
    .C(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__a21oi_1 _18074_ (.A1(_02353_),
    .A2(_02354_),
    .B1(_02355_),
    .Y(_02357_));
 sky130_fd_sc_hd__o31a_1 _18075_ (.A1(_02341_),
    .A2(_02356_),
    .A3(_02357_),
    .B1(_02337_),
    .X(_02358_));
 sky130_fd_sc_hd__o2bb2a_1 _18076_ (.A1_N(_09830_),
    .A2_N(_02358_),
    .B1(_02340_),
    .B2(\rbzero.wall_tracer.trackDistY[-8] ),
    .X(_00553_));
 sky130_fd_sc_hd__nor2_1 _18077_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_02359_));
 sky130_fd_sc_hd__nand2_1 _18078_ (.A(\rbzero.wall_tracer.trackDistY[-7] ),
    .B(\rbzero.wall_tracer.stepDistY[-7] ),
    .Y(_02360_));
 sky130_fd_sc_hd__or2b_1 _18079_ (.A(_02359_),
    .B_N(_02360_),
    .X(_02361_));
 sky130_fd_sc_hd__a21boi_1 _18080_ (.A1(_02353_),
    .A2(_02355_),
    .B1_N(_02354_),
    .Y(_02362_));
 sky130_fd_sc_hd__xnor2_1 _18081_ (.A(_02361_),
    .B(_02362_),
    .Y(_02363_));
 sky130_fd_sc_hd__clkbuf_4 _18082_ (.A(_02336_),
    .X(_02364_));
 sky130_fd_sc_hd__o21a_1 _18083_ (.A1(_09872_),
    .A2(_02363_),
    .B1(_02364_),
    .X(_02365_));
 sky130_fd_sc_hd__o2bb2a_1 _18084_ (.A1_N(_09837_),
    .A2_N(_02365_),
    .B1(_02340_),
    .B2(\rbzero.wall_tracer.trackDistY[-7] ),
    .X(_00554_));
 sky130_fd_sc_hd__or2_1 _18085_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .X(_02366_));
 sky130_fd_sc_hd__nand2_1 _18086_ (.A(\rbzero.wall_tracer.trackDistY[-6] ),
    .B(\rbzero.wall_tracer.stepDistY[-6] ),
    .Y(_02367_));
 sky130_fd_sc_hd__o21ai_1 _18087_ (.A1(_02359_),
    .A2(_02362_),
    .B1(_02360_),
    .Y(_02368_));
 sky130_fd_sc_hd__a21oi_1 _18088_ (.A1(_02366_),
    .A2(_02367_),
    .B1(_02368_),
    .Y(_02369_));
 sky130_fd_sc_hd__a31o_1 _18089_ (.A1(_02366_),
    .A2(_02367_),
    .A3(_02368_),
    .B1(_06104_),
    .X(_02370_));
 sky130_fd_sc_hd__o21a_1 _18090_ (.A1(_02369_),
    .A2(_02370_),
    .B1(_02364_),
    .X(_02371_));
 sky130_fd_sc_hd__o2bb2a_1 _18091_ (.A1_N(_09845_),
    .A2_N(_02371_),
    .B1(_02340_),
    .B2(\rbzero.wall_tracer.trackDistY[-6] ),
    .X(_00555_));
 sky130_fd_sc_hd__nor2_1 _18092_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_02372_));
 sky130_fd_sc_hd__nand2_1 _18093_ (.A(\rbzero.wall_tracer.trackDistY[-5] ),
    .B(\rbzero.wall_tracer.stepDistY[-5] ),
    .Y(_02373_));
 sky130_fd_sc_hd__or2b_1 _18094_ (.A(_02372_),
    .B_N(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__a21boi_1 _18095_ (.A1(_02366_),
    .A2(_02368_),
    .B1_N(_02367_),
    .Y(_02375_));
 sky130_fd_sc_hd__nor2_1 _18096_ (.A(_02374_),
    .B(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__a21o_1 _18097_ (.A1(_02374_),
    .A2(_02375_),
    .B1(_09866_),
    .X(_02377_));
 sky130_fd_sc_hd__o21ai_1 _18098_ (.A1(_02376_),
    .A2(_02377_),
    .B1(_09852_),
    .Y(_02378_));
 sky130_fd_sc_hd__mux2_1 _18099_ (.A0(\rbzero.wall_tracer.trackDistY[-5] ),
    .A1(_02378_),
    .S(_02339_),
    .X(_02379_));
 sky130_fd_sc_hd__clkbuf_1 _18100_ (.A(_02379_),
    .X(_00556_));
 sky130_fd_sc_hd__or2_1 _18101_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .X(_02380_));
 sky130_fd_sc_hd__nand2_1 _18102_ (.A(\rbzero.wall_tracer.trackDistY[-4] ),
    .B(\rbzero.wall_tracer.stepDistY[-4] ),
    .Y(_02381_));
 sky130_fd_sc_hd__o21ai_1 _18103_ (.A1(_02372_),
    .A2(_02375_),
    .B1(_02373_),
    .Y(_02382_));
 sky130_fd_sc_hd__a21oi_1 _18104_ (.A1(_02380_),
    .A2(_02381_),
    .B1(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__a31o_1 _18105_ (.A1(_02380_),
    .A2(_02381_),
    .A3(_02382_),
    .B1(_06104_),
    .X(_02384_));
 sky130_fd_sc_hd__o21a_1 _18106_ (.A1(_02383_),
    .A2(_02384_),
    .B1(_02337_),
    .X(_02385_));
 sky130_fd_sc_hd__o2bb2a_1 _18107_ (.A1_N(_09859_),
    .A2_N(_02385_),
    .B1(_02340_),
    .B2(\rbzero.wall_tracer.trackDistY[-4] ),
    .X(_00557_));
 sky130_fd_sc_hd__nor2_1 _18108_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_02386_));
 sky130_fd_sc_hd__nand2_1 _18109_ (.A(\rbzero.wall_tracer.trackDistY[-3] ),
    .B(\rbzero.wall_tracer.stepDistY[-3] ),
    .Y(_02387_));
 sky130_fd_sc_hd__or2b_1 _18110_ (.A(_02386_),
    .B_N(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__a21boi_1 _18111_ (.A1(_02380_),
    .A2(_02382_),
    .B1_N(_02381_),
    .Y(_02389_));
 sky130_fd_sc_hd__nor2_1 _18112_ (.A(_02388_),
    .B(_02389_),
    .Y(_02390_));
 sky130_fd_sc_hd__a21o_1 _18113_ (.A1(_02388_),
    .A2(_02389_),
    .B1(_09866_),
    .X(_02391_));
 sky130_fd_sc_hd__o21ai_1 _18114_ (.A1(_02390_),
    .A2(_02391_),
    .B1(_09869_),
    .Y(_02392_));
 sky130_fd_sc_hd__mux2_1 _18115_ (.A0(\rbzero.wall_tracer.trackDistY[-3] ),
    .A1(_02392_),
    .S(_02339_),
    .X(_02393_));
 sky130_fd_sc_hd__clkbuf_1 _18116_ (.A(_02393_),
    .X(_00558_));
 sky130_fd_sc_hd__or2_1 _18117_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .X(_02394_));
 sky130_fd_sc_hd__nand2_1 _18118_ (.A(\rbzero.wall_tracer.trackDistY[-2] ),
    .B(\rbzero.wall_tracer.stepDistY[-2] ),
    .Y(_02395_));
 sky130_fd_sc_hd__o21ai_1 _18119_ (.A1(_02386_),
    .A2(_02389_),
    .B1(_02387_),
    .Y(_02396_));
 sky130_fd_sc_hd__and3_1 _18120_ (.A(_02394_),
    .B(_02395_),
    .C(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__a21oi_1 _18121_ (.A1(_02394_),
    .A2(_02395_),
    .B1(_02396_),
    .Y(_02398_));
 sky130_fd_sc_hd__o31a_1 _18122_ (.A1(_02341_),
    .A2(_02397_),
    .A3(_02398_),
    .B1(_02337_),
    .X(_02399_));
 sky130_fd_sc_hd__o2bb2a_1 _18123_ (.A1_N(_09873_),
    .A2_N(_02399_),
    .B1(_02340_),
    .B2(\rbzero.wall_tracer.trackDistY[-2] ),
    .X(_00559_));
 sky130_fd_sc_hd__nor2_1 _18124_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .Y(_02400_));
 sky130_fd_sc_hd__and2_1 _18125_ (.A(\rbzero.wall_tracer.trackDistY[-1] ),
    .B(\rbzero.wall_tracer.stepDistY[-1] ),
    .X(_02401_));
 sky130_fd_sc_hd__a21boi_1 _18126_ (.A1(_02394_),
    .A2(_02396_),
    .B1_N(_02395_),
    .Y(_02402_));
 sky130_fd_sc_hd__nor3_1 _18127_ (.A(_02400_),
    .B(_02401_),
    .C(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__o21a_1 _18128_ (.A1(_02400_),
    .A2(_02401_),
    .B1(_02402_),
    .X(_02404_));
 sky130_fd_sc_hd__o31a_1 _18129_ (.A1(_02341_),
    .A2(_02403_),
    .A3(_02404_),
    .B1(_02339_),
    .X(_02405_));
 sky130_fd_sc_hd__o2bb2a_1 _18130_ (.A1_N(_09887_),
    .A2_N(_02405_),
    .B1(_02340_),
    .B2(\rbzero.wall_tracer.trackDistY[-1] ),
    .X(_00560_));
 sky130_fd_sc_hd__or2_1 _18131_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .X(_02406_));
 sky130_fd_sc_hd__nand2_1 _18132_ (.A(\rbzero.wall_tracer.trackDistY[0] ),
    .B(\rbzero.wall_tracer.stepDistY[0] ),
    .Y(_02407_));
 sky130_fd_sc_hd__a211oi_1 _18133_ (.A1(_02406_),
    .A2(_02407_),
    .B1(_02401_),
    .C1(_02403_),
    .Y(_02408_));
 sky130_fd_sc_hd__o211a_1 _18134_ (.A1(_02401_),
    .A2(_02403_),
    .B1(_02406_),
    .C1(_02407_),
    .X(_02409_));
 sky130_fd_sc_hd__o31a_1 _18135_ (.A1(_02341_),
    .A2(_02408_),
    .A3(_02409_),
    .B1(_02339_),
    .X(_02410_));
 sky130_fd_sc_hd__o2bb2a_1 _18136_ (.A1_N(_10011_),
    .A2_N(_02410_),
    .B1(_02340_),
    .B2(\rbzero.wall_tracer.trackDistY[0] ),
    .X(_00561_));
 sky130_fd_sc_hd__nand2_1 _18137_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .Y(_02411_));
 sky130_fd_sc_hd__or2_1 _18138_ (.A(\rbzero.wall_tracer.trackDistY[1] ),
    .B(\rbzero.wall_tracer.stepDistY[1] ),
    .X(_02412_));
 sky130_fd_sc_hd__a21o_1 _18139_ (.A1(\rbzero.wall_tracer.trackDistY[0] ),
    .A2(\rbzero.wall_tracer.stepDistY[0] ),
    .B1(_02409_),
    .X(_02413_));
 sky130_fd_sc_hd__and3_1 _18140_ (.A(_02411_),
    .B(_02412_),
    .C(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__a21oi_1 _18141_ (.A1(_02411_),
    .A2(_02412_),
    .B1(_02413_),
    .Y(_02415_));
 sky130_fd_sc_hd__o31a_1 _18142_ (.A1(_02341_),
    .A2(_02414_),
    .A3(_02415_),
    .B1(_02339_),
    .X(_02416_));
 sky130_fd_sc_hd__o2bb2a_1 _18143_ (.A1_N(_10127_),
    .A2_N(_02416_),
    .B1(_02364_),
    .B2(\rbzero.wall_tracer.trackDistY[1] ),
    .X(_00562_));
 sky130_fd_sc_hd__nand2_1 _18144_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .Y(_02417_));
 sky130_fd_sc_hd__or2_1 _18145_ (.A(\rbzero.wall_tracer.trackDistY[2] ),
    .B(\rbzero.wall_tracer.stepDistY[2] ),
    .X(_02418_));
 sky130_fd_sc_hd__inv_2 _18146_ (.A(_02411_),
    .Y(_02419_));
 sky130_fd_sc_hd__a211o_1 _18147_ (.A1(_02417_),
    .A2(_02418_),
    .B1(_02419_),
    .C1(_02414_),
    .X(_02420_));
 sky130_fd_sc_hd__o211ai_2 _18148_ (.A1(_02419_),
    .A2(_02414_),
    .B1(_02417_),
    .C1(_02418_),
    .Y(_02421_));
 sky130_fd_sc_hd__nand2_1 _18149_ (.A(_02420_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__o21a_1 _18150_ (.A1(_09872_),
    .A2(_02422_),
    .B1(_02337_),
    .X(_02423_));
 sky130_fd_sc_hd__o2bb2a_1 _18151_ (.A1_N(_10259_),
    .A2_N(_02423_),
    .B1(_02364_),
    .B2(\rbzero.wall_tracer.trackDistY[2] ),
    .X(_00563_));
 sky130_fd_sc_hd__and2_1 _18152_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .X(_02424_));
 sky130_fd_sc_hd__nor2_1 _18153_ (.A(\rbzero.wall_tracer.trackDistY[3] ),
    .B(\rbzero.wall_tracer.stepDistY[3] ),
    .Y(_02425_));
 sky130_fd_sc_hd__o211a_1 _18154_ (.A1(_02424_),
    .A2(_02425_),
    .B1(_02417_),
    .C1(_02421_),
    .X(_02426_));
 sky130_fd_sc_hd__a211oi_2 _18155_ (.A1(_02417_),
    .A2(_02421_),
    .B1(_02424_),
    .C1(_02425_),
    .Y(_02427_));
 sky130_fd_sc_hd__o31a_1 _18156_ (.A1(_02341_),
    .A2(_02426_),
    .A3(_02427_),
    .B1(_02339_),
    .X(_02428_));
 sky130_fd_sc_hd__o2bb2a_1 _18157_ (.A1_N(_10375_),
    .A2_N(_02428_),
    .B1(_02364_),
    .B2(\rbzero.wall_tracer.trackDistY[3] ),
    .X(_00564_));
 sky130_fd_sc_hd__nand2_1 _18158_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .Y(_02429_));
 sky130_fd_sc_hd__or2_1 _18159_ (.A(\rbzero.wall_tracer.trackDistY[4] ),
    .B(\rbzero.wall_tracer.stepDistY[4] ),
    .X(_02430_));
 sky130_fd_sc_hd__o211a_1 _18160_ (.A1(_02424_),
    .A2(_02427_),
    .B1(_02429_),
    .C1(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__a211oi_1 _18161_ (.A1(_02429_),
    .A2(_02430_),
    .B1(_02424_),
    .C1(_02427_),
    .Y(_02432_));
 sky130_fd_sc_hd__o31a_1 _18162_ (.A1(_02341_),
    .A2(_02431_),
    .A3(_02432_),
    .B1(_02339_),
    .X(_02433_));
 sky130_fd_sc_hd__o2bb2a_1 _18163_ (.A1_N(_01759_),
    .A2_N(_02433_),
    .B1(_02364_),
    .B2(\rbzero.wall_tracer.trackDistY[4] ),
    .X(_00565_));
 sky130_fd_sc_hd__nor2_1 _18164_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .Y(_02434_));
 sky130_fd_sc_hd__and2_1 _18165_ (.A(\rbzero.wall_tracer.trackDistY[5] ),
    .B(\rbzero.wall_tracer.stepDistY[5] ),
    .X(_02435_));
 sky130_fd_sc_hd__a21oi_1 _18166_ (.A1(\rbzero.wall_tracer.trackDistY[4] ),
    .A2(\rbzero.wall_tracer.stepDistY[4] ),
    .B1(_02431_),
    .Y(_02436_));
 sky130_fd_sc_hd__nor3_1 _18167_ (.A(_02434_),
    .B(_02435_),
    .C(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__o21a_1 _18168_ (.A1(_02434_),
    .A2(_02435_),
    .B1(_02436_),
    .X(_02438_));
 sky130_fd_sc_hd__o31a_1 _18169_ (.A1(_02341_),
    .A2(_02437_),
    .A3(_02438_),
    .B1(_02339_),
    .X(_02439_));
 sky130_fd_sc_hd__o2bb2a_1 _18170_ (.A1_N(_01868_),
    .A2_N(_02439_),
    .B1(_02364_),
    .B2(\rbzero.wall_tracer.trackDistY[5] ),
    .X(_00566_));
 sky130_fd_sc_hd__nor2_1 _18171_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .Y(_02440_));
 sky130_fd_sc_hd__and2_1 _18172_ (.A(\rbzero.wall_tracer.trackDistY[6] ),
    .B(\rbzero.wall_tracer.stepDistY[6] ),
    .X(_02441_));
 sky130_fd_sc_hd__o21ba_1 _18173_ (.A1(_02434_),
    .A2(_02436_),
    .B1_N(_02435_),
    .X(_02442_));
 sky130_fd_sc_hd__o21ai_1 _18174_ (.A1(_02440_),
    .A2(_02441_),
    .B1(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__o31a_1 _18175_ (.A1(_02440_),
    .A2(_02441_),
    .A3(_02442_),
    .B1(_08123_),
    .X(_02444_));
 sky130_fd_sc_hd__a21bo_1 _18176_ (.A1(_02443_),
    .A2(_02444_),
    .B1_N(_01981_),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _18177_ (.A0(\rbzero.wall_tracer.trackDistY[6] ),
    .A1(_02445_),
    .S(_02339_),
    .X(_02446_));
 sky130_fd_sc_hd__clkbuf_1 _18178_ (.A(_02446_),
    .X(_00567_));
 sky130_fd_sc_hd__nor2_1 _18179_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_02447_));
 sky130_fd_sc_hd__nand2_1 _18180_ (.A(\rbzero.wall_tracer.trackDistY[7] ),
    .B(\rbzero.wall_tracer.stepDistY[7] ),
    .Y(_02448_));
 sky130_fd_sc_hd__or2b_1 _18181_ (.A(_02447_),
    .B_N(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__o21ba_1 _18182_ (.A1(_02440_),
    .A2(_02442_),
    .B1_N(_02441_),
    .X(_02450_));
 sky130_fd_sc_hd__nor2_1 _18183_ (.A(_02449_),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__a21o_1 _18184_ (.A1(_02449_),
    .A2(_02450_),
    .B1(_09866_),
    .X(_02452_));
 sky130_fd_sc_hd__o21ai_1 _18185_ (.A1(_02451_),
    .A2(_02452_),
    .B1(_02083_),
    .Y(_02453_));
 sky130_fd_sc_hd__mux2_1 _18186_ (.A0(\rbzero.wall_tracer.trackDistY[7] ),
    .A1(_02453_),
    .S(_02336_),
    .X(_02454_));
 sky130_fd_sc_hd__clkbuf_1 _18187_ (.A(_02454_),
    .X(_00568_));
 sky130_fd_sc_hd__or2_1 _18188_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .X(_02455_));
 sky130_fd_sc_hd__nand2_1 _18189_ (.A(\rbzero.wall_tracer.trackDistY[8] ),
    .B(\rbzero.wall_tracer.stepDistY[8] ),
    .Y(_02456_));
 sky130_fd_sc_hd__nand2_1 _18190_ (.A(_02455_),
    .B(_02456_),
    .Y(_02457_));
 sky130_fd_sc_hd__o21a_1 _18191_ (.A1(_02447_),
    .A2(_02450_),
    .B1(_02448_),
    .X(_02458_));
 sky130_fd_sc_hd__nor2_1 _18192_ (.A(_02457_),
    .B(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__a21o_1 _18193_ (.A1(_02457_),
    .A2(_02458_),
    .B1(_06104_),
    .X(_02460_));
 sky130_fd_sc_hd__o21a_1 _18194_ (.A1(_02459_),
    .A2(_02460_),
    .B1(_02337_),
    .X(_02461_));
 sky130_fd_sc_hd__o2bb2a_1 _18195_ (.A1_N(_02176_),
    .A2_N(_02461_),
    .B1(_02364_),
    .B2(\rbzero.wall_tracer.trackDistY[8] ),
    .X(_00569_));
 sky130_fd_sc_hd__and2_1 _18196_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .X(_02462_));
 sky130_fd_sc_hd__nor2_1 _18197_ (.A(\rbzero.wall_tracer.trackDistY[9] ),
    .B(\rbzero.wall_tracer.stepDistY[9] ),
    .Y(_02463_));
 sky130_fd_sc_hd__nor2_1 _18198_ (.A(_02462_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2_1 _18199_ (.A(_02456_),
    .B(_02458_),
    .Y(_02465_));
 sky130_fd_sc_hd__and2_1 _18200_ (.A(_02455_),
    .B(_02465_),
    .X(_02466_));
 sky130_fd_sc_hd__xnor2_1 _18201_ (.A(_02464_),
    .B(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__o21a_1 _18202_ (.A1(_09872_),
    .A2(_02467_),
    .B1(_02337_),
    .X(_02468_));
 sky130_fd_sc_hd__o2bb2a_1 _18203_ (.A1_N(_02262_),
    .A2_N(_02468_),
    .B1(_02364_),
    .B2(\rbzero.wall_tracer.trackDistY[9] ),
    .X(_00570_));
 sky130_fd_sc_hd__a31o_1 _18204_ (.A1(_02455_),
    .A2(_02464_),
    .A3(_02465_),
    .B1(_02462_),
    .X(_02469_));
 sky130_fd_sc_hd__xor2_1 _18205_ (.A(\rbzero.wall_tracer.trackDistY[10] ),
    .B(\rbzero.wall_tracer.stepDistY[10] ),
    .X(_02470_));
 sky130_fd_sc_hd__xnor2_1 _18206_ (.A(_02469_),
    .B(_02470_),
    .Y(_02471_));
 sky130_fd_sc_hd__o21a_1 _18207_ (.A1(_09872_),
    .A2(_02471_),
    .B1(_02337_),
    .X(_02472_));
 sky130_fd_sc_hd__o2bb2a_1 _18208_ (.A1_N(_02329_),
    .A2_N(_02472_),
    .B1(_02364_),
    .B2(\rbzero.wall_tracer.trackDistY[10] ),
    .X(_00571_));
 sky130_fd_sc_hd__buf_4 _18209_ (.A(\rbzero.spi_registers.spi_buffer[0] ),
    .X(_02473_));
 sky130_fd_sc_hd__buf_2 _18210_ (.A(\rbzero.spi_registers.spi_cmd[1] ),
    .X(_02474_));
 sky130_fd_sc_hd__clkbuf_2 _18211_ (.A(\rbzero.spi_registers.spi_cmd[2] ),
    .X(_02475_));
 sky130_fd_sc_hd__inv_2 _18212_ (.A(\rbzero.spi_registers.spi_cmd[3] ),
    .Y(_02476_));
 sky130_fd_sc_hd__or4b_4 _18213_ (.A(_02475_),
    .B(_02476_),
    .C(_04052_),
    .D_N(\rbzero.spi_registers.spi_done ),
    .X(_02477_));
 sky130_fd_sc_hd__nor3b_4 _18214_ (.A(_02474_),
    .B(_02477_),
    .C_N(\rbzero.spi_registers.spi_cmd[0] ),
    .Y(_02478_));
 sky130_fd_sc_hd__buf_4 _18215_ (.A(_02478_),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _18216_ (.A0(\rbzero.spi_registers.new_texadd[2][0] ),
    .A1(_02473_),
    .S(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__clkbuf_1 _18217_ (.A(_02480_),
    .X(_00572_));
 sky130_fd_sc_hd__buf_4 _18218_ (.A(\rbzero.spi_registers.spi_buffer[1] ),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _18219_ (.A0(\rbzero.spi_registers.new_texadd[2][1] ),
    .A1(_02481_),
    .S(_02479_),
    .X(_02482_));
 sky130_fd_sc_hd__clkbuf_1 _18220_ (.A(_02482_),
    .X(_00573_));
 sky130_fd_sc_hd__buf_4 _18221_ (.A(\rbzero.spi_registers.spi_buffer[2] ),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _18222_ (.A0(\rbzero.spi_registers.new_texadd[2][2] ),
    .A1(_02483_),
    .S(_02479_),
    .X(_02484_));
 sky130_fd_sc_hd__clkbuf_1 _18223_ (.A(_02484_),
    .X(_00574_));
 sky130_fd_sc_hd__buf_4 _18224_ (.A(\rbzero.spi_registers.spi_buffer[3] ),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _18225_ (.A0(\rbzero.spi_registers.new_texadd[2][3] ),
    .A1(_02485_),
    .S(_02479_),
    .X(_02486_));
 sky130_fd_sc_hd__clkbuf_1 _18226_ (.A(_02486_),
    .X(_00575_));
 sky130_fd_sc_hd__buf_4 _18227_ (.A(\rbzero.spi_registers.spi_buffer[4] ),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _18228_ (.A0(\rbzero.spi_registers.new_texadd[2][4] ),
    .A1(_02487_),
    .S(_02479_),
    .X(_02488_));
 sky130_fd_sc_hd__clkbuf_1 _18229_ (.A(_02488_),
    .X(_00576_));
 sky130_fd_sc_hd__clkbuf_4 _18230_ (.A(\rbzero.spi_registers.spi_buffer[5] ),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _18231_ (.A0(\rbzero.spi_registers.new_texadd[2][5] ),
    .A1(_02489_),
    .S(_02479_),
    .X(_02490_));
 sky130_fd_sc_hd__clkbuf_1 _18232_ (.A(_02490_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _18233_ (.A0(\rbzero.spi_registers.new_texadd[2][6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_02479_),
    .X(_02491_));
 sky130_fd_sc_hd__clkbuf_1 _18234_ (.A(_02491_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _18235_ (.A0(\rbzero.spi_registers.new_texadd[2][7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_02479_),
    .X(_02492_));
 sky130_fd_sc_hd__clkbuf_1 _18236_ (.A(_02492_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _18237_ (.A0(\rbzero.spi_registers.new_texadd[2][8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_02479_),
    .X(_02493_));
 sky130_fd_sc_hd__clkbuf_1 _18238_ (.A(_02493_),
    .X(_00580_));
 sky130_fd_sc_hd__buf_4 _18239_ (.A(_02478_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _18240_ (.A0(\rbzero.spi_registers.new_texadd[2][9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__clkbuf_1 _18241_ (.A(_02495_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _18242_ (.A0(\rbzero.spi_registers.new_texadd[2][10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_02494_),
    .X(_02496_));
 sky130_fd_sc_hd__clkbuf_1 _18243_ (.A(_02496_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _18244_ (.A0(\rbzero.spi_registers.new_texadd[2][11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_02494_),
    .X(_02497_));
 sky130_fd_sc_hd__clkbuf_1 _18245_ (.A(_02497_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _18246_ (.A0(\rbzero.spi_registers.new_texadd[2][12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_02494_),
    .X(_02498_));
 sky130_fd_sc_hd__clkbuf_1 _18247_ (.A(_02498_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _18248_ (.A0(\rbzero.spi_registers.new_texadd[2][13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_02494_),
    .X(_02499_));
 sky130_fd_sc_hd__clkbuf_1 _18249_ (.A(_02499_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _18250_ (.A0(\rbzero.spi_registers.new_texadd[2][14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_02494_),
    .X(_02500_));
 sky130_fd_sc_hd__clkbuf_1 _18251_ (.A(_02500_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _18252_ (.A0(\rbzero.spi_registers.new_texadd[2][15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_02494_),
    .X(_02501_));
 sky130_fd_sc_hd__clkbuf_1 _18253_ (.A(_02501_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _18254_ (.A0(\rbzero.spi_registers.new_texadd[2][16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_02494_),
    .X(_02502_));
 sky130_fd_sc_hd__clkbuf_1 _18255_ (.A(_02502_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _18256_ (.A0(\rbzero.spi_registers.new_texadd[2][17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_02494_),
    .X(_02503_));
 sky130_fd_sc_hd__clkbuf_1 _18257_ (.A(_02503_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _18258_ (.A0(\rbzero.spi_registers.new_texadd[2][18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_02494_),
    .X(_02504_));
 sky130_fd_sc_hd__clkbuf_1 _18259_ (.A(_02504_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _18260_ (.A0(\rbzero.spi_registers.new_texadd[2][19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_02478_),
    .X(_02505_));
 sky130_fd_sc_hd__clkbuf_1 _18261_ (.A(_02505_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _18262_ (.A0(\rbzero.spi_registers.new_texadd[2][20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_02478_),
    .X(_02506_));
 sky130_fd_sc_hd__clkbuf_1 _18263_ (.A(_02506_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _18264_ (.A0(\rbzero.spi_registers.new_texadd[2][21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_02478_),
    .X(_02507_));
 sky130_fd_sc_hd__clkbuf_1 _18265_ (.A(_02507_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _18266_ (.A0(\rbzero.spi_registers.new_texadd[2][22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_02478_),
    .X(_02508_));
 sky130_fd_sc_hd__clkbuf_1 _18267_ (.A(_02508_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _18268_ (.A0(\rbzero.spi_registers.new_texadd[2][23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_02478_),
    .X(_02509_));
 sky130_fd_sc_hd__clkbuf_1 _18269_ (.A(_02509_),
    .X(_00595_));
 sky130_fd_sc_hd__nor2_1 _18270_ (.A(_05111_),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_02510_));
 sky130_fd_sc_hd__nand2_1 _18271_ (.A(_05111_),
    .B(\rbzero.wall_tracer.rayAddendX[-5] ),
    .Y(_02511_));
 sky130_fd_sc_hd__and2b_1 _18272_ (.A_N(_02510_),
    .B(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__nor2_1 _18273_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_02513_));
 sky130_fd_sc_hd__nand2_1 _18274_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .Y(_02514_));
 sky130_fd_sc_hd__nor2_1 _18275_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .Y(_02515_));
 sky130_fd_sc_hd__and2_1 _18276_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.wall_tracer.rayAddendX[-8] ),
    .X(_02516_));
 sky130_fd_sc_hd__o21ba_1 _18277_ (.A1(_02514_),
    .A2(_02515_),
    .B1_N(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__nand2_1 _18278_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(\rbzero.wall_tracer.rayAddendX[-7] ),
    .Y(_02518_));
 sky130_fd_sc_hd__o21ai_1 _18279_ (.A1(_02513_),
    .A2(_02517_),
    .B1(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__a21o_1 _18280_ (.A1(\rbzero.debug_overlay.vplaneX[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[-6] ),
    .B1(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__o21ai_1 _18281_ (.A1(_05120_),
    .A2(\rbzero.wall_tracer.rayAddendX[-6] ),
    .B1(_02520_),
    .Y(_02521_));
 sky130_fd_sc_hd__xnor2_1 _18282_ (.A(_02512_),
    .B(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__mux2_1 _18283_ (.A0(\rbzero.debug_overlay.vplaneX[-9] ),
    .A1(_02522_),
    .S(_04433_),
    .X(_02523_));
 sky130_fd_sc_hd__or2_1 _18284_ (.A(_04432_),
    .B(_09743_),
    .X(_02524_));
 sky130_fd_sc_hd__buf_4 _18285_ (.A(_02524_),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _18286_ (.A0(\rbzero.wall_tracer.rayAddendX[-5] ),
    .A1(_02523_),
    .S(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__clkbuf_1 _18287_ (.A(_02526_),
    .X(_00596_));
 sky130_fd_sc_hd__buf_4 _18288_ (.A(_02525_),
    .X(_02527_));
 sky130_fd_sc_hd__nor2_1 _18289_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .Y(_02528_));
 sky130_fd_sc_hd__and2_1 _18290_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(_02529_));
 sky130_fd_sc_hd__o21ai_1 _18291_ (.A1(_02510_),
    .A2(_02521_),
    .B1(_02511_),
    .Y(_02530_));
 sky130_fd_sc_hd__or3_1 _18292_ (.A(_02528_),
    .B(_02529_),
    .C(_02530_),
    .X(_02531_));
 sky130_fd_sc_hd__o21ai_1 _18293_ (.A1(_02528_),
    .A2(_02529_),
    .B1(_02530_),
    .Y(_02532_));
 sky130_fd_sc_hd__a21oi_1 _18294_ (.A1(_02531_),
    .A2(_02532_),
    .B1(_08136_),
    .Y(_02533_));
 sky130_fd_sc_hd__clkbuf_4 _18295_ (.A(_08135_),
    .X(_02534_));
 sky130_fd_sc_hd__nand2_1 _18296_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .Y(_02535_));
 sky130_fd_sc_hd__or2_1 _18297_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(\rbzero.debug_overlay.vplaneX[-9] ),
    .X(_02536_));
 sky130_fd_sc_hd__a31o_1 _18298_ (.A1(_02534_),
    .A2(_02535_),
    .A3(_02536_),
    .B1(_09745_),
    .X(_02537_));
 sky130_fd_sc_hd__o22a_1 _18299_ (.A1(\rbzero.wall_tracer.rayAddendX[-4] ),
    .A2(_02527_),
    .B1(_02533_),
    .B2(_02537_),
    .X(_00597_));
 sky130_fd_sc_hd__nor2_1 _18300_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02538_));
 sky130_fd_sc_hd__and2_1 _18301_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .X(_02539_));
 sky130_fd_sc_hd__or2_1 _18302_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.wall_tracer.rayAddendX[-4] ),
    .X(_02540_));
 sky130_fd_sc_hd__a21oi_1 _18303_ (.A1(_02540_),
    .A2(_02530_),
    .B1(_02529_),
    .Y(_02541_));
 sky130_fd_sc_hd__o21ai_1 _18304_ (.A1(_02538_),
    .A2(_02539_),
    .B1(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__o311a_1 _18305_ (.A1(_02538_),
    .A2(_02539_),
    .A3(_02541_),
    .B1(_02542_),
    .C1(_04442_),
    .X(_02543_));
 sky130_fd_sc_hd__or2_1 _18306_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_02536_),
    .X(_02544_));
 sky130_fd_sc_hd__nand2_1 _18307_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_02536_),
    .Y(_02545_));
 sky130_fd_sc_hd__a31o_1 _18308_ (.A1(_02534_),
    .A2(_02544_),
    .A3(_02545_),
    .B1(_09745_),
    .X(_02546_));
 sky130_fd_sc_hd__o22a_1 _18309_ (.A1(\rbzero.wall_tracer.rayAddendX[-3] ),
    .A2(_02527_),
    .B1(_02543_),
    .B2(_02546_),
    .X(_00598_));
 sky130_fd_sc_hd__nor2_1 _18310_ (.A(_05106_),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .Y(_02547_));
 sky130_fd_sc_hd__and2_1 _18311_ (.A(_05106_),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_02548_));
 sky130_fd_sc_hd__nand2_1 _18312_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.wall_tracer.rayAddendX[-3] ),
    .Y(_02549_));
 sky130_fd_sc_hd__o21ai_1 _18313_ (.A1(_02538_),
    .A2(_02541_),
    .B1(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__or3_1 _18314_ (.A(_02547_),
    .B(_02548_),
    .C(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__o21ai_1 _18315_ (.A1(_02547_),
    .A2(_02548_),
    .B1(_02550_),
    .Y(_02552_));
 sky130_fd_sc_hd__a21oi_1 _18316_ (.A1(_02551_),
    .A2(_02552_),
    .B1(_08136_),
    .Y(_02553_));
 sky130_fd_sc_hd__nand2_1 _18317_ (.A(_05120_),
    .B(_02544_),
    .Y(_02554_));
 sky130_fd_sc_hd__or2_1 _18318_ (.A(_05120_),
    .B(_02544_),
    .X(_02555_));
 sky130_fd_sc_hd__a31o_1 _18319_ (.A1(_02534_),
    .A2(_02554_),
    .A3(_02555_),
    .B1(_09745_),
    .X(_02556_));
 sky130_fd_sc_hd__o22a_1 _18320_ (.A1(\rbzero.wall_tracer.rayAddendX[-2] ),
    .A2(_02527_),
    .B1(_02553_),
    .B2(_02556_),
    .X(_00599_));
 sky130_fd_sc_hd__buf_6 _18321_ (.A(_09749_),
    .X(_02557_));
 sky130_fd_sc_hd__or2_1 _18322_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .X(_02558_));
 sky130_fd_sc_hd__nand2_1 _18323_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(\rbzero.wall_tracer.rayAddendX[-1] ),
    .Y(_02559_));
 sky130_fd_sc_hd__or2_1 _18324_ (.A(\rbzero.debug_overlay.vplaneX[-2] ),
    .B(\rbzero.wall_tracer.rayAddendX[-2] ),
    .X(_02560_));
 sky130_fd_sc_hd__a21o_1 _18325_ (.A1(_02560_),
    .A2(_02550_),
    .B1(_02548_),
    .X(_02561_));
 sky130_fd_sc_hd__nand3_1 _18326_ (.A(_02558_),
    .B(_02559_),
    .C(_02561_),
    .Y(_02562_));
 sky130_fd_sc_hd__a21o_1 _18327_ (.A1(_02558_),
    .A2(_02559_),
    .B1(_02561_),
    .X(_02563_));
 sky130_fd_sc_hd__inv_2 _18328_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .Y(_02564_));
 sky130_fd_sc_hd__o31a_1 _18329_ (.A1(_05120_),
    .A2(\rbzero.debug_overlay.vplaneX[-7] ),
    .A3(\rbzero.debug_overlay.vplaneX[-8] ),
    .B1(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__xor2_1 _18330_ (.A(_05111_),
    .B(_02565_),
    .X(_02566_));
 sky130_fd_sc_hd__a22o_1 _18331_ (.A1(\rbzero.wall_tracer.rayAddendX[-1] ),
    .A2(_09745_),
    .B1(_02566_),
    .B2(_02534_),
    .X(_02567_));
 sky130_fd_sc_hd__a31o_1 _18332_ (.A1(_02557_),
    .A2(_02562_),
    .A3(_02563_),
    .B1(_02567_),
    .X(_00600_));
 sky130_fd_sc_hd__a21bo_1 _18333_ (.A1(_02558_),
    .A2(_02561_),
    .B1_N(_02559_),
    .X(_02568_));
 sky130_fd_sc_hd__clkbuf_4 _18334_ (.A(\rbzero.debug_overlay.vplaneX[0] ),
    .X(_02569_));
 sky130_fd_sc_hd__nor2_1 _18335_ (.A(_02569_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .Y(_02570_));
 sky130_fd_sc_hd__and2_1 _18336_ (.A(_02569_),
    .B(\rbzero.wall_tracer.rayAddendX[0] ),
    .X(_02571_));
 sky130_fd_sc_hd__or2_1 _18337_ (.A(_02570_),
    .B(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__xnor2_1 _18338_ (.A(_02568_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__or2_1 _18339_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .X(_02574_));
 sky130_fd_sc_hd__nand2_1 _18340_ (.A(\rbzero.debug_overlay.vplaneX[-4] ),
    .B(\rbzero.debug_overlay.vplaneX[-8] ),
    .Y(_02575_));
 sky130_fd_sc_hd__nand2_1 _18341_ (.A(_02574_),
    .B(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__nor2_1 _18342_ (.A(_05111_),
    .B(_02555_),
    .Y(_02577_));
 sky130_fd_sc_hd__a21oi_1 _18343_ (.A1(_05111_),
    .A2(\rbzero.debug_overlay.vplaneX[-9] ),
    .B1(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__xnor2_1 _18344_ (.A(_02576_),
    .B(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__mux2_1 _18345_ (.A0(_02573_),
    .A1(_02579_),
    .S(_08134_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _18346_ (.A0(\rbzero.wall_tracer.rayAddendX[0] ),
    .A1(_02580_),
    .S(_02525_),
    .X(_02581_));
 sky130_fd_sc_hd__clkbuf_1 _18347_ (.A(_02581_),
    .X(_00601_));
 sky130_fd_sc_hd__nand2_1 _18348_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .Y(_02582_));
 sky130_fd_sc_hd__or2_1 _18349_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .B(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02583_));
 sky130_fd_sc_hd__o21a_1 _18350_ (.A1(_02569_),
    .A2(\rbzero.wall_tracer.rayAddendX[0] ),
    .B1(_02568_),
    .X(_02584_));
 sky130_fd_sc_hd__a211o_1 _18351_ (.A1(_02582_),
    .A2(_02583_),
    .B1(_02584_),
    .C1(_02571_),
    .X(_02585_));
 sky130_fd_sc_hd__o211ai_2 _18352_ (.A1(_02571_),
    .A2(_02584_),
    .B1(_02583_),
    .C1(_02582_),
    .Y(_02586_));
 sky130_fd_sc_hd__a21oi_1 _18353_ (.A1(_05111_),
    .A2(\rbzero.debug_overlay.vplaneX[-9] ),
    .B1(_02576_),
    .Y(_02587_));
 sky130_fd_sc_hd__nor2_1 _18354_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .Y(_02588_));
 sky130_fd_sc_hd__and2_1 _18355_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(\rbzero.debug_overlay.vplaneX[-7] ),
    .X(_02589_));
 sky130_fd_sc_hd__nor2_1 _18356_ (.A(_02588_),
    .B(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__xnor2_1 _18357_ (.A(_02574_),
    .B(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__o21a_1 _18358_ (.A1(_02577_),
    .A2(_02587_),
    .B1(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__inv_2 _18359_ (.A(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__or3_1 _18360_ (.A(_02577_),
    .B(_02591_),
    .C(_02587_),
    .X(_02594_));
 sky130_fd_sc_hd__a32o_1 _18361_ (.A1(_08135_),
    .A2(_02593_),
    .A3(_02594_),
    .B1(_09751_),
    .B2(\rbzero.wall_tracer.rayAddendX[1] ),
    .X(_02595_));
 sky130_fd_sc_hd__a31o_1 _18362_ (.A1(_02557_),
    .A2(_02585_),
    .A3(_02586_),
    .B1(_02595_),
    .X(_00602_));
 sky130_fd_sc_hd__buf_2 _18363_ (.A(\rbzero.debug_overlay.vplaneX[10] ),
    .X(_02596_));
 sky130_fd_sc_hd__buf_2 _18364_ (.A(_02596_),
    .X(_02597_));
 sky130_fd_sc_hd__clkbuf_4 _18365_ (.A(_02597_),
    .X(_02598_));
 sky130_fd_sc_hd__xnor2_1 _18366_ (.A(_02598_),
    .B(\rbzero.wall_tracer.rayAddendX[2] ),
    .Y(_02599_));
 sky130_fd_sc_hd__a21oi_1 _18367_ (.A1(_02582_),
    .A2(_02586_),
    .B1(_02599_),
    .Y(_02600_));
 sky130_fd_sc_hd__a311oi_1 _18368_ (.A1(_02582_),
    .A2(_02586_),
    .A3(_02599_),
    .B1(_02600_),
    .C1(_08136_),
    .Y(_02601_));
 sky130_fd_sc_hd__xor2_1 _18369_ (.A(_05106_),
    .B(_05120_),
    .X(_02602_));
 sky130_fd_sc_hd__o31ai_1 _18370_ (.A1(_02574_),
    .A2(_02588_),
    .A3(_02589_),
    .B1(_02593_),
    .Y(_02603_));
 sky130_fd_sc_hd__xnor2_1 _18371_ (.A(_02602_),
    .B(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__xnor2_1 _18372_ (.A(_02588_),
    .B(_02604_),
    .Y(_02605_));
 sky130_fd_sc_hd__buf_6 _18373_ (.A(_09744_),
    .X(_02606_));
 sky130_fd_sc_hd__a21o_1 _18374_ (.A1(_08136_),
    .A2(_02605_),
    .B1(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__o22a_1 _18375_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(_02527_),
    .B1(_02601_),
    .B2(_02607_),
    .X(_00603_));
 sky130_fd_sc_hd__and2_1 _18376_ (.A(_02596_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .X(_02608_));
 sky130_fd_sc_hd__nor2_1 _18377_ (.A(_02596_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02609_));
 sky130_fd_sc_hd__o21ai_1 _18378_ (.A1(\rbzero.wall_tracer.rayAddendX[2] ),
    .A2(\rbzero.wall_tracer.rayAddendX[1] ),
    .B1(_02596_),
    .Y(_02610_));
 sky130_fd_sc_hd__o21bai_1 _18379_ (.A1(_02596_),
    .A2(\rbzero.wall_tracer.rayAddendX[2] ),
    .B1_N(_02586_),
    .Y(_02611_));
 sky130_fd_sc_hd__o211ai_1 _18380_ (.A1(_02608_),
    .A2(_02609_),
    .B1(_02610_),
    .C1(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__a211o_1 _18381_ (.A1(_02610_),
    .A2(_02611_),
    .B1(_02608_),
    .C1(_02609_),
    .X(_02613_));
 sky130_fd_sc_hd__or2_1 _18382_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_05111_),
    .X(_02614_));
 sky130_fd_sc_hd__nand2_1 _18383_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_05111_),
    .Y(_02615_));
 sky130_fd_sc_hd__and4bb_1 _18384_ (.A_N(_05106_),
    .B_N(_05120_),
    .C(_02614_),
    .D(_02615_),
    .X(_02616_));
 sky130_fd_sc_hd__a2bb2o_1 _18385_ (.A1_N(_05106_),
    .A2_N(_05120_),
    .B1(_02614_),
    .B2(_02615_),
    .X(_02617_));
 sky130_fd_sc_hd__and2b_1 _18386_ (.A_N(_02616_),
    .B(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__o21a_1 _18387_ (.A1(_02592_),
    .A2(_02602_),
    .B1(_02588_),
    .X(_02619_));
 sky130_fd_sc_hd__a21o_1 _18388_ (.A1(_02602_),
    .A2(_02603_),
    .B1(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__and2_1 _18389_ (.A(_02618_),
    .B(_02620_),
    .X(_02621_));
 sky130_fd_sc_hd__o21ai_1 _18390_ (.A1(_02618_),
    .A2(_02620_),
    .B1(_08135_),
    .Y(_02622_));
 sky130_fd_sc_hd__a2bb2o_1 _18391_ (.A1_N(_02621_),
    .A2_N(_02622_),
    .B1(\rbzero.wall_tracer.rayAddendX[3] ),
    .B2(_09744_),
    .X(_02623_));
 sky130_fd_sc_hd__a31o_1 _18392_ (.A1(_02557_),
    .A2(_02612_),
    .A3(_02613_),
    .B1(_02623_),
    .X(_00604_));
 sky130_fd_sc_hd__nand2_1 _18393_ (.A(_02598_),
    .B(\rbzero.wall_tracer.rayAddendX[3] ),
    .Y(_02624_));
 sky130_fd_sc_hd__xor2_1 _18394_ (.A(_02596_),
    .B(\rbzero.wall_tracer.rayAddendX[4] ),
    .X(_02625_));
 sky130_fd_sc_hd__a21oi_1 _18395_ (.A1(_02624_),
    .A2(_02613_),
    .B1(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hd__a31o_1 _18396_ (.A1(_02624_),
    .A2(_02613_),
    .A3(_02625_),
    .B1(_08134_),
    .X(_02627_));
 sky130_fd_sc_hd__xor2_1 _18397_ (.A(_02569_),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .X(_02628_));
 sky130_fd_sc_hd__o21ai_1 _18398_ (.A1(_02616_),
    .A2(_02621_),
    .B1(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hd__or3_1 _18399_ (.A(_02616_),
    .B(_02621_),
    .C(_02628_),
    .X(_02630_));
 sky130_fd_sc_hd__and2_1 _18400_ (.A(_02629_),
    .B(_02630_),
    .X(_02631_));
 sky130_fd_sc_hd__xnor2_1 _18401_ (.A(_02614_),
    .B(_02631_),
    .Y(_02632_));
 sky130_fd_sc_hd__o22a_1 _18402_ (.A1(_02626_),
    .A2(_02627_),
    .B1(_02632_),
    .B2(_04434_),
    .X(_02633_));
 sky130_fd_sc_hd__mux2_1 _18403_ (.A0(\rbzero.wall_tracer.rayAddendX[4] ),
    .A1(_02633_),
    .S(_02525_),
    .X(_02634_));
 sky130_fd_sc_hd__clkbuf_1 _18404_ (.A(_02634_),
    .X(_00605_));
 sky130_fd_sc_hd__nand2_1 _18405_ (.A(_02597_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .Y(_02635_));
 sky130_fd_sc_hd__or2_1 _18406_ (.A(_02596_),
    .B(\rbzero.wall_tracer.rayAddendX[5] ),
    .X(_02636_));
 sky130_fd_sc_hd__nand2_1 _18407_ (.A(_02635_),
    .B(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hd__or2b_1 _18408_ (.A(_02613_),
    .B_N(_02625_),
    .X(_02638_));
 sky130_fd_sc_hd__o21ai_1 _18409_ (.A1(\rbzero.wall_tracer.rayAddendX[4] ),
    .A2(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02598_),
    .Y(_02639_));
 sky130_fd_sc_hd__nand3_1 _18410_ (.A(_02637_),
    .B(_02638_),
    .C(_02639_),
    .Y(_02640_));
 sky130_fd_sc_hd__a21o_1 _18411_ (.A1(_02638_),
    .A2(_02639_),
    .B1(_02637_),
    .X(_02641_));
 sky130_fd_sc_hd__nor2_1 _18412_ (.A(_02596_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .Y(_02642_));
 sky130_fd_sc_hd__and2_1 _18413_ (.A(_02596_),
    .B(\rbzero.debug_overlay.vplaneX[-3] ),
    .X(_02643_));
 sky130_fd_sc_hd__o22a_1 _18414_ (.A1(_02569_),
    .A2(\rbzero.debug_overlay.vplaneX[-4] ),
    .B1(_02642_),
    .B2(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__nor4_1 _18415_ (.A(_02569_),
    .B(\rbzero.debug_overlay.vplaneX[-4] ),
    .C(_02642_),
    .D(_02643_),
    .Y(_02645_));
 sky130_fd_sc_hd__nor2_1 _18416_ (.A(_02644_),
    .B(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__a2bb2o_1 _18417_ (.A1_N(_02621_),
    .A2_N(_02628_),
    .B1(_02629_),
    .B2(_02614_),
    .X(_02647_));
 sky130_fd_sc_hd__xnor2_1 _18418_ (.A(_02646_),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__a22o_1 _18419_ (.A1(\rbzero.wall_tracer.rayAddendX[5] ),
    .A2(_09745_),
    .B1(_02648_),
    .B2(_02534_),
    .X(_02649_));
 sky130_fd_sc_hd__a31o_1 _18420_ (.A1(_09753_),
    .A2(_02640_),
    .A3(_02641_),
    .B1(_02649_),
    .X(_00606_));
 sky130_fd_sc_hd__xnor2_1 _18421_ (.A(_02597_),
    .B(\rbzero.wall_tracer.rayAddendX[6] ),
    .Y(_02650_));
 sky130_fd_sc_hd__a21oi_1 _18422_ (.A1(_02635_),
    .A2(_02641_),
    .B1(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hd__a31o_1 _18423_ (.A1(_02635_),
    .A2(_02641_),
    .A3(_02650_),
    .B1(_08134_),
    .X(_02652_));
 sky130_fd_sc_hd__or2_1 _18424_ (.A(_02596_),
    .B(_05106_),
    .X(_02653_));
 sky130_fd_sc_hd__nand2_1 _18425_ (.A(_02597_),
    .B(_05106_),
    .Y(_02654_));
 sky130_fd_sc_hd__a21o_1 _18426_ (.A1(_02653_),
    .A2(_02654_),
    .B1(_02642_),
    .X(_02655_));
 sky130_fd_sc_hd__nand2_1 _18427_ (.A(_05106_),
    .B(_02642_),
    .Y(_02656_));
 sky130_fd_sc_hd__nand2_1 _18428_ (.A(_02655_),
    .B(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__o21bai_1 _18429_ (.A1(_02644_),
    .A2(_02647_),
    .B1_N(_02645_),
    .Y(_02658_));
 sky130_fd_sc_hd__xnor2_1 _18430_ (.A(_02657_),
    .B(_02658_),
    .Y(_02659_));
 sky130_fd_sc_hd__a2bb2o_1 _18431_ (.A1_N(_02651_),
    .A2_N(_02652_),
    .B1(_02659_),
    .B2(_08134_),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _18432_ (.A0(\rbzero.wall_tracer.rayAddendX[6] ),
    .A1(_02660_),
    .S(_02525_),
    .X(_02661_));
 sky130_fd_sc_hd__clkbuf_1 _18433_ (.A(_02661_),
    .X(_00607_));
 sky130_fd_sc_hd__nand2_1 _18434_ (.A(_02597_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .Y(_02662_));
 sky130_fd_sc_hd__or2_1 _18435_ (.A(_02597_),
    .B(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02663_));
 sky130_fd_sc_hd__nor3_1 _18436_ (.A(_02637_),
    .B(_02638_),
    .C(_02650_),
    .Y(_02664_));
 sky130_fd_sc_hd__o41a_1 _18437_ (.A1(\rbzero.wall_tracer.rayAddendX[6] ),
    .A2(\rbzero.wall_tracer.rayAddendX[5] ),
    .A3(\rbzero.wall_tracer.rayAddendX[4] ),
    .A4(\rbzero.wall_tracer.rayAddendX[3] ),
    .B1(_02597_),
    .X(_02665_));
 sky130_fd_sc_hd__a211o_1 _18438_ (.A1(_02662_),
    .A2(_02663_),
    .B1(_02664_),
    .C1(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__o211ai_2 _18439_ (.A1(_02664_),
    .A2(_02665_),
    .B1(_02662_),
    .C1(_02663_),
    .Y(_02667_));
 sky130_fd_sc_hd__inv_2 _18440_ (.A(_02656_),
    .Y(_02668_));
 sky130_fd_sc_hd__and3_1 _18441_ (.A(_02655_),
    .B(_02656_),
    .C(_02658_),
    .X(_02669_));
 sky130_fd_sc_hd__nor2_1 _18442_ (.A(_02597_),
    .B(\rbzero.debug_overlay.vplaneX[-1] ),
    .Y(_02670_));
 sky130_fd_sc_hd__and2_1 _18443_ (.A(_02597_),
    .B(\rbzero.debug_overlay.vplaneX[-1] ),
    .X(_02671_));
 sky130_fd_sc_hd__o21ai_1 _18444_ (.A1(_02670_),
    .A2(_02671_),
    .B1(_02653_),
    .Y(_02672_));
 sky130_fd_sc_hd__or3_1 _18445_ (.A(_02653_),
    .B(_02670_),
    .C(_02671_),
    .X(_02673_));
 sky130_fd_sc_hd__o211ai_2 _18446_ (.A1(_02668_),
    .A2(_02669_),
    .B1(_02672_),
    .C1(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__a211o_1 _18447_ (.A1(_02672_),
    .A2(_02673_),
    .B1(_02668_),
    .C1(_02669_),
    .X(_02675_));
 sky130_fd_sc_hd__a32o_1 _18448_ (.A1(_08135_),
    .A2(_02674_),
    .A3(_02675_),
    .B1(_09751_),
    .B2(\rbzero.wall_tracer.rayAddendX[7] ),
    .X(_02676_));
 sky130_fd_sc_hd__a31o_1 _18449_ (.A1(_09753_),
    .A2(_02666_),
    .A3(_02667_),
    .B1(_02676_),
    .X(_00608_));
 sky130_fd_sc_hd__xnor2_1 _18450_ (.A(_02597_),
    .B(\rbzero.wall_tracer.rayAddendX[8] ),
    .Y(_02677_));
 sky130_fd_sc_hd__a21oi_1 _18451_ (.A1(_02662_),
    .A2(_02667_),
    .B1(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__a31o_1 _18452_ (.A1(_02662_),
    .A2(_02667_),
    .A3(_02677_),
    .B1(_08135_),
    .X(_02679_));
 sky130_fd_sc_hd__nor2_1 _18453_ (.A(_02678_),
    .B(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__inv_2 _18454_ (.A(_02569_),
    .Y(_02681_));
 sky130_fd_sc_hd__a21oi_1 _18455_ (.A1(_02569_),
    .A2(\rbzero.debug_overlay.vplaneX[-1] ),
    .B1(_02598_),
    .Y(_02682_));
 sky130_fd_sc_hd__a21oi_1 _18456_ (.A1(_02598_),
    .A2(_02569_),
    .B1(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__a21oi_1 _18457_ (.A1(_02681_),
    .A2(_02670_),
    .B1(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__a21o_1 _18458_ (.A1(_02673_),
    .A2(_02674_),
    .B1(_02684_),
    .X(_02685_));
 sky130_fd_sc_hd__nand3_1 _18459_ (.A(_02673_),
    .B(_02674_),
    .C(_02684_),
    .Y(_02686_));
 sky130_fd_sc_hd__a31o_1 _18460_ (.A1(_02534_),
    .A2(_02685_),
    .A3(_02686_),
    .B1(_09745_),
    .X(_02687_));
 sky130_fd_sc_hd__o22a_1 _18461_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(_02527_),
    .B1(_02680_),
    .B2(_02687_),
    .X(_00609_));
 sky130_fd_sc_hd__or2_1 _18462_ (.A(_02598_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .X(_02688_));
 sky130_fd_sc_hd__nand2_1 _18463_ (.A(_02598_),
    .B(\rbzero.wall_tracer.rayAddendX[9] ),
    .Y(_02689_));
 sky130_fd_sc_hd__nand2_1 _18464_ (.A(_02688_),
    .B(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__o21ai_1 _18465_ (.A1(\rbzero.wall_tracer.rayAddendX[8] ),
    .A2(\rbzero.wall_tracer.rayAddendX[7] ),
    .B1(_02598_),
    .Y(_02691_));
 sky130_fd_sc_hd__o21ai_1 _18466_ (.A1(_02667_),
    .A2(_02677_),
    .B1(_02691_),
    .Y(_02692_));
 sky130_fd_sc_hd__xnor2_1 _18467_ (.A(_02690_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__inv_2 _18468_ (.A(_02598_),
    .Y(_02694_));
 sky130_fd_sc_hd__a21oi_1 _18469_ (.A1(_02694_),
    .A2(_02681_),
    .B1(_02685_),
    .Y(_02695_));
 sky130_fd_sc_hd__a211o_1 _18470_ (.A1(_02682_),
    .A2(_02685_),
    .B1(_02695_),
    .C1(_04434_),
    .X(_02696_));
 sky130_fd_sc_hd__o221a_1 _18471_ (.A1(\rbzero.wall_tracer.rayAddendX[9] ),
    .A2(_02527_),
    .B1(_09760_),
    .B2(_02693_),
    .C1(_02696_),
    .X(_00610_));
 sky130_fd_sc_hd__a21bo_1 _18472_ (.A1(_02688_),
    .A2(_02692_),
    .B1_N(_02689_),
    .X(_02697_));
 sky130_fd_sc_hd__xnor2_1 _18473_ (.A(_02598_),
    .B(\rbzero.wall_tracer.rayAddendX[10] ),
    .Y(_02698_));
 sky130_fd_sc_hd__xnor2_1 _18474_ (.A(_02697_),
    .B(_02698_),
    .Y(_02699_));
 sky130_fd_sc_hd__o21a_1 _18475_ (.A1(_02569_),
    .A2(_02685_),
    .B1(_08134_),
    .X(_02700_));
 sky130_fd_sc_hd__a22o_1 _18476_ (.A1(_04434_),
    .A2(_02699_),
    .B1(_02700_),
    .B2(_02694_),
    .X(_02701_));
 sky130_fd_sc_hd__mux2_1 _18477_ (.A0(\rbzero.wall_tracer.rayAddendX[10] ),
    .A1(_02701_),
    .S(_02525_),
    .X(_02702_));
 sky130_fd_sc_hd__clkbuf_1 _18478_ (.A(_02702_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _18479_ (.A0(\rbzero.debug_overlay.playerY[0] ),
    .A1(_06130_),
    .S(_01757_),
    .X(_02703_));
 sky130_fd_sc_hd__o21a_2 _18480_ (.A1(_06161_),
    .A2(_06258_),
    .B1(_06264_),
    .X(_02704_));
 sky130_fd_sc_hd__mux2_1 _18481_ (.A0(_06088_),
    .A1(_02703_),
    .S(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__clkbuf_1 _18482_ (.A(_02705_),
    .X(_00612_));
 sky130_fd_sc_hd__nor2_1 _18483_ (.A(_06088_),
    .B(_06090_),
    .Y(_02706_));
 sky130_fd_sc_hd__or3_1 _18484_ (.A(_09866_),
    .B(_06091_),
    .C(_02706_),
    .X(_02707_));
 sky130_fd_sc_hd__o211a_1 _18485_ (.A1(_06111_),
    .A2(_08124_),
    .B1(_02704_),
    .C1(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__a21oi_1 _18486_ (.A1(_06089_),
    .A2(_06265_),
    .B1(_02708_),
    .Y(_00613_));
 sky130_fd_sc_hd__nor2_1 _18487_ (.A(_06092_),
    .B(_06093_),
    .Y(_02709_));
 sky130_fd_sc_hd__nand2_1 _18488_ (.A(_08124_),
    .B(_06094_),
    .Y(_02710_));
 sky130_fd_sc_hd__o221a_1 _18489_ (.A1(_06112_),
    .A2(_08124_),
    .B1(_02709_),
    .B2(_02710_),
    .C1(_02704_),
    .X(_02711_));
 sky130_fd_sc_hd__a21oi_1 _18490_ (.A1(_06086_),
    .A2(_06265_),
    .B1(_02711_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_1 _18491_ (.A(_06084_),
    .B(_06096_),
    .Y(_02712_));
 sky130_fd_sc_hd__xnor2_1 _18492_ (.A(_06095_),
    .B(_02712_),
    .Y(_02713_));
 sky130_fd_sc_hd__mux2_1 _18493_ (.A0(\rbzero.debug_overlay.playerY[3] ),
    .A1(_02713_),
    .S(_01757_),
    .X(_02714_));
 sky130_fd_sc_hd__mux2_1 _18494_ (.A0(\rbzero.map_rom.a6 ),
    .A1(_02714_),
    .S(_02704_),
    .X(_02715_));
 sky130_fd_sc_hd__clkbuf_1 _18495_ (.A(_02715_),
    .X(_00615_));
 sky130_fd_sc_hd__nand2_1 _18496_ (.A(_06082_),
    .B(_06083_),
    .Y(_02716_));
 sky130_fd_sc_hd__xnor2_1 _18497_ (.A(_02716_),
    .B(_06097_),
    .Y(_02717_));
 sky130_fd_sc_hd__mux2_1 _18498_ (.A0(\rbzero.debug_overlay.playerY[4] ),
    .A1(_02717_),
    .S(_01757_),
    .X(_02718_));
 sky130_fd_sc_hd__mux2_1 _18499_ (.A0(\rbzero.map_rom.i_row[4] ),
    .A1(_02718_),
    .S(_02704_),
    .X(_02719_));
 sky130_fd_sc_hd__clkbuf_1 _18500_ (.A(_02719_),
    .X(_00616_));
 sky130_fd_sc_hd__a21oi_1 _18501_ (.A1(\rbzero.map_rom.i_row[4] ),
    .A2(_06078_),
    .B1(_06098_),
    .Y(_02720_));
 sky130_fd_sc_hd__xnor2_1 _18502_ (.A(_06081_),
    .B(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__mux2_1 _18503_ (.A0(\rbzero.debug_overlay.playerY[5] ),
    .A1(_02721_),
    .S(_01757_),
    .X(_02722_));
 sky130_fd_sc_hd__mux2_1 _18504_ (.A0(\rbzero.wall_tracer.mapY[5] ),
    .A1(_02722_),
    .S(_02704_),
    .X(_02723_));
 sky130_fd_sc_hd__clkbuf_1 _18505_ (.A(_02723_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _18506_ (.A0(\rbzero.debug_overlay.playerX[0] ),
    .A1(_06108_),
    .S(_01757_),
    .X(_02724_));
 sky130_fd_sc_hd__mux2_1 _18507_ (.A0(_06144_),
    .A1(_02724_),
    .S(_09844_),
    .X(_02725_));
 sky130_fd_sc_hd__clkbuf_1 _18508_ (.A(_02725_),
    .X(_00618_));
 sky130_fd_sc_hd__nor2_1 _18509_ (.A(_06144_),
    .B(_09766_),
    .Y(_02726_));
 sky130_fd_sc_hd__or3_1 _18510_ (.A(_09866_),
    .B(_09767_),
    .C(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__o211a_1 _18511_ (.A1(_04671_),
    .A2(_08124_),
    .B1(_09844_),
    .C1(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__a21oi_1 _18512_ (.A1(_06117_),
    .A2(_09785_),
    .B1(_02728_),
    .Y(_00619_));
 sky130_fd_sc_hd__xnor2_1 _18513_ (.A(_09768_),
    .B(_09771_),
    .Y(_02729_));
 sky130_fd_sc_hd__mux2_1 _18514_ (.A0(_04674_),
    .A1(_02729_),
    .S(_08124_),
    .X(_02730_));
 sky130_fd_sc_hd__nor2_1 _18515_ (.A(\rbzero.map_rom.f2 ),
    .B(_09879_),
    .Y(_02731_));
 sky130_fd_sc_hd__a21oi_1 _18516_ (.A1(_09879_),
    .A2(_02730_),
    .B1(_02731_),
    .Y(_00620_));
 sky130_fd_sc_hd__or2b_1 _18517_ (.A(_09765_),
    .B_N(_09773_),
    .X(_02732_));
 sky130_fd_sc_hd__xnor2_1 _18518_ (.A(_09772_),
    .B(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__mux2_1 _18519_ (.A0(\rbzero.debug_overlay.playerX[3] ),
    .A1(_02733_),
    .S(_01757_),
    .X(_02734_));
 sky130_fd_sc_hd__mux2_1 _18520_ (.A0(\rbzero.map_rom.f1 ),
    .A1(_02734_),
    .S(_09844_),
    .X(_02735_));
 sky130_fd_sc_hd__clkbuf_1 _18521_ (.A(_02735_),
    .X(_00621_));
 sky130_fd_sc_hd__xnor2_1 _18522_ (.A(_09775_),
    .B(_09774_),
    .Y(_02736_));
 sky130_fd_sc_hd__mux2_1 _18523_ (.A0(\rbzero.debug_overlay.playerX[4] ),
    .A1(_02736_),
    .S(_01757_),
    .X(_02737_));
 sky130_fd_sc_hd__mux2_1 _18524_ (.A0(\rbzero.map_rom.i_col[4] ),
    .A1(_02737_),
    .S(_09844_),
    .X(_02738_));
 sky130_fd_sc_hd__clkbuf_1 _18525_ (.A(_02738_),
    .X(_00622_));
 sky130_fd_sc_hd__a21oi_1 _18526_ (.A1(\rbzero.map_rom.i_col[4] ),
    .A2(_09119_),
    .B1(_09776_),
    .Y(_02739_));
 sky130_fd_sc_hd__xnor2_1 _18527_ (.A(_09764_),
    .B(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__mux2_1 _18528_ (.A0(\rbzero.debug_overlay.playerX[5] ),
    .A1(_02740_),
    .S(_08123_),
    .X(_02741_));
 sky130_fd_sc_hd__mux2_1 _18529_ (.A0(\rbzero.wall_tracer.mapX[5] ),
    .A1(_02741_),
    .S(_09844_),
    .X(_02742_));
 sky130_fd_sc_hd__clkbuf_1 _18530_ (.A(_02742_),
    .X(_00623_));
 sky130_fd_sc_hd__nor2_1 _18531_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_02743_));
 sky130_fd_sc_hd__nand2_1 _18532_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.wall_tracer.rayAddendY[-5] ),
    .Y(_02744_));
 sky130_fd_sc_hd__and2b_1 _18533_ (.A_N(_02743_),
    .B(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__nor2_1 _18534_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_02746_));
 sky130_fd_sc_hd__nand2_1 _18535_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .Y(_02747_));
 sky130_fd_sc_hd__nor2_1 _18536_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .Y(_02748_));
 sky130_fd_sc_hd__and2_1 _18537_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.wall_tracer.rayAddendY[-8] ),
    .X(_02749_));
 sky130_fd_sc_hd__o21ba_1 _18538_ (.A1(_02747_),
    .A2(_02748_),
    .B1_N(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__nand2_1 _18539_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(\rbzero.wall_tracer.rayAddendY[-7] ),
    .Y(_02751_));
 sky130_fd_sc_hd__o21ai_1 _18540_ (.A1(_02746_),
    .A2(_02750_),
    .B1(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__a21o_1 _18541_ (.A1(\rbzero.debug_overlay.vplaneY[-6] ),
    .A2(\rbzero.wall_tracer.rayAddendY[-6] ),
    .B1(_02752_),
    .X(_02753_));
 sky130_fd_sc_hd__o21ai_1 _18542_ (.A1(_05129_),
    .A2(\rbzero.wall_tracer.rayAddendY[-6] ),
    .B1(_02753_),
    .Y(_02754_));
 sky130_fd_sc_hd__xnor2_1 _18543_ (.A(_02745_),
    .B(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__inv_2 _18544_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_02756_));
 sky130_fd_sc_hd__nor2_1 _18545_ (.A(_02756_),
    .B(_04442_),
    .Y(_02757_));
 sky130_fd_sc_hd__a221o_1 _18546_ (.A1(\rbzero.wall_tracer.rayAddendY[-5] ),
    .A2(_02606_),
    .B1(_09753_),
    .B2(_02755_),
    .C1(_02757_),
    .X(_00624_));
 sky130_fd_sc_hd__nor2_1 _18547_ (.A(_05132_),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .Y(_02758_));
 sky130_fd_sc_hd__and2_1 _18548_ (.A(_05132_),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_02759_));
 sky130_fd_sc_hd__o21ai_1 _18549_ (.A1(_02743_),
    .A2(_02754_),
    .B1(_02744_),
    .Y(_02760_));
 sky130_fd_sc_hd__or3_1 _18550_ (.A(_02758_),
    .B(_02759_),
    .C(_02760_),
    .X(_02761_));
 sky130_fd_sc_hd__o21ai_1 _18551_ (.A1(_02758_),
    .A2(_02759_),
    .B1(_02760_),
    .Y(_02762_));
 sky130_fd_sc_hd__a21oi_1 _18552_ (.A1(_02761_),
    .A2(_02762_),
    .B1(_08136_),
    .Y(_02763_));
 sky130_fd_sc_hd__or2_1 _18553_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .X(_02764_));
 sky130_fd_sc_hd__nand2_1 _18554_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_02765_));
 sky130_fd_sc_hd__a31o_1 _18555_ (.A1(_02534_),
    .A2(_02764_),
    .A3(_02765_),
    .B1(_09745_),
    .X(_02766_));
 sky130_fd_sc_hd__o22a_1 _18556_ (.A1(\rbzero.wall_tracer.rayAddendY[-4] ),
    .A2(_02527_),
    .B1(_02763_),
    .B2(_02766_),
    .X(_00625_));
 sky130_fd_sc_hd__nor2_1 _18557_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02767_));
 sky130_fd_sc_hd__and2_1 _18558_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .X(_02768_));
 sky130_fd_sc_hd__or2_1 _18559_ (.A(\rbzero.debug_overlay.vplaneY[-4] ),
    .B(\rbzero.wall_tracer.rayAddendY[-4] ),
    .X(_02769_));
 sky130_fd_sc_hd__a21oi_1 _18560_ (.A1(_02769_),
    .A2(_02760_),
    .B1(_02759_),
    .Y(_02770_));
 sky130_fd_sc_hd__o21ai_1 _18561_ (.A1(_02767_),
    .A2(_02768_),
    .B1(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__o311a_1 _18562_ (.A1(_02767_),
    .A2(_02768_),
    .A3(_02770_),
    .B1(_02771_),
    .C1(_04442_),
    .X(_02772_));
 sky130_fd_sc_hd__or2_1 _18563_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_02764_),
    .X(_02773_));
 sky130_fd_sc_hd__nand2_1 _18564_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_02764_),
    .Y(_02774_));
 sky130_fd_sc_hd__a31o_1 _18565_ (.A1(_08135_),
    .A2(_02773_),
    .A3(_02774_),
    .B1(_09745_),
    .X(_02775_));
 sky130_fd_sc_hd__o22a_1 _18566_ (.A1(\rbzero.wall_tracer.rayAddendY[-3] ),
    .A2(_02527_),
    .B1(_02772_),
    .B2(_02775_),
    .X(_00626_));
 sky130_fd_sc_hd__or2_1 _18567_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .X(_02776_));
 sky130_fd_sc_hd__nand2_1 _18568_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(\rbzero.wall_tracer.rayAddendY[-2] ),
    .Y(_02777_));
 sky130_fd_sc_hd__nand2_1 _18569_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.wall_tracer.rayAddendY[-3] ),
    .Y(_02778_));
 sky130_fd_sc_hd__o21ai_1 _18570_ (.A1(_02767_),
    .A2(_02770_),
    .B1(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__a21oi_1 _18571_ (.A1(_02776_),
    .A2(_02777_),
    .B1(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__a31o_1 _18572_ (.A1(_02776_),
    .A2(_02777_),
    .A3(_02779_),
    .B1(_08134_),
    .X(_02781_));
 sky130_fd_sc_hd__or2_1 _18573_ (.A(_05129_),
    .B(_02773_),
    .X(_02782_));
 sky130_fd_sc_hd__a21oi_1 _18574_ (.A1(_05129_),
    .A2(_02773_),
    .B1(_04433_),
    .Y(_02783_));
 sky130_fd_sc_hd__a2bb2o_1 _18575_ (.A1_N(_02780_),
    .A2_N(_02781_),
    .B1(_02782_),
    .B2(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__mux2_1 _18576_ (.A0(\rbzero.wall_tracer.rayAddendY[-2] ),
    .A1(_02784_),
    .S(_02525_),
    .X(_02785_));
 sky130_fd_sc_hd__clkbuf_1 _18577_ (.A(_02785_),
    .X(_00627_));
 sky130_fd_sc_hd__or2_1 _18578_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .X(_02786_));
 sky130_fd_sc_hd__nand2_1 _18579_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.wall_tracer.rayAddendY[-1] ),
    .Y(_02787_));
 sky130_fd_sc_hd__a21bo_1 _18580_ (.A1(_02776_),
    .A2(_02779_),
    .B1_N(_02777_),
    .X(_02788_));
 sky130_fd_sc_hd__nand3_1 _18581_ (.A(_02786_),
    .B(_02787_),
    .C(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__a21o_1 _18582_ (.A1(_02786_),
    .A2(_02787_),
    .B1(_02788_),
    .X(_02790_));
 sky130_fd_sc_hd__o31a_1 _18583_ (.A1(_05129_),
    .A2(\rbzero.debug_overlay.vplaneY[-7] ),
    .A3(\rbzero.debug_overlay.vplaneY[-8] ),
    .B1(_02756_),
    .X(_02791_));
 sky130_fd_sc_hd__xor2_1 _18584_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__a22o_1 _18585_ (.A1(\rbzero.wall_tracer.rayAddendY[-1] ),
    .A2(_09744_),
    .B1(_02792_),
    .B2(_02534_),
    .X(_02793_));
 sky130_fd_sc_hd__a31o_1 _18586_ (.A1(_09753_),
    .A2(_02789_),
    .A3(_02790_),
    .B1(_02793_),
    .X(_00628_));
 sky130_fd_sc_hd__clkbuf_4 _18587_ (.A(\rbzero.debug_overlay.vplaneY[0] ),
    .X(_02794_));
 sky130_fd_sc_hd__nor2_1 _18588_ (.A(_02794_),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .Y(_02795_));
 sky130_fd_sc_hd__and2_1 _18589_ (.A(_02794_),
    .B(\rbzero.wall_tracer.rayAddendY[0] ),
    .X(_02796_));
 sky130_fd_sc_hd__a21bo_1 _18590_ (.A1(_02786_),
    .A2(_02788_),
    .B1_N(_02787_),
    .X(_02797_));
 sky130_fd_sc_hd__o21ai_1 _18591_ (.A1(_02795_),
    .A2(_02796_),
    .B1(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__o31a_1 _18592_ (.A1(_02797_),
    .A2(_02795_),
    .A3(_02796_),
    .B1(_04433_),
    .X(_02799_));
 sky130_fd_sc_hd__or2_1 _18593_ (.A(_05132_),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .X(_02800_));
 sky130_fd_sc_hd__nand2_1 _18594_ (.A(_05132_),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .Y(_02801_));
 sky130_fd_sc_hd__nand2_1 _18595_ (.A(_02800_),
    .B(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_1 _18596_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(\rbzero.debug_overlay.vplaneY[-9] ),
    .Y(_02803_));
 sky130_fd_sc_hd__or2_1 _18597_ (.A(\rbzero.debug_overlay.vplaneY[-5] ),
    .B(_02782_),
    .X(_02804_));
 sky130_fd_sc_hd__nand2_1 _18598_ (.A(_02803_),
    .B(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__xor2_1 _18599_ (.A(_02802_),
    .B(_02805_),
    .X(_02806_));
 sky130_fd_sc_hd__o2bb2a_1 _18600_ (.A1_N(_02798_),
    .A2_N(_02799_),
    .B1(_02806_),
    .B2(_04434_),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _18601_ (.A0(\rbzero.wall_tracer.rayAddendY[0] ),
    .A1(_02807_),
    .S(_02525_),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_1 _18602_ (.A(_02808_),
    .X(_00629_));
 sky130_fd_sc_hd__nand2_1 _18603_ (.A(_05127_),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .Y(_02809_));
 sky130_fd_sc_hd__or2_1 _18604_ (.A(\rbzero.debug_overlay.vplaneY[10] ),
    .B(\rbzero.wall_tracer.rayAddendY[1] ),
    .X(_02810_));
 sky130_fd_sc_hd__o21a_1 _18605_ (.A1(_02794_),
    .A2(\rbzero.wall_tracer.rayAddendY[0] ),
    .B1(_02797_),
    .X(_02811_));
 sky130_fd_sc_hd__a211o_1 _18606_ (.A1(_02809_),
    .A2(_02810_),
    .B1(_02811_),
    .C1(_02796_),
    .X(_02812_));
 sky130_fd_sc_hd__o211ai_2 _18607_ (.A1(_02796_),
    .A2(_02811_),
    .B1(_02810_),
    .C1(_02809_),
    .Y(_02813_));
 sky130_fd_sc_hd__nor2_1 _18608_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .Y(_02814_));
 sky130_fd_sc_hd__and2_1 _18609_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(\rbzero.debug_overlay.vplaneY[-7] ),
    .X(_02815_));
 sky130_fd_sc_hd__nor2_1 _18610_ (.A(_02814_),
    .B(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__xnor2_1 _18611_ (.A(_02800_),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__a21bo_1 _18612_ (.A1(_02802_),
    .A2(_02804_),
    .B1_N(_02803_),
    .X(_02818_));
 sky130_fd_sc_hd__xnor2_1 _18613_ (.A(_02817_),
    .B(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__a22o_1 _18614_ (.A1(\rbzero.wall_tracer.rayAddendY[1] ),
    .A2(_09744_),
    .B1(_02819_),
    .B2(_02534_),
    .X(_02820_));
 sky130_fd_sc_hd__a31o_1 _18615_ (.A1(_09753_),
    .A2(_02812_),
    .A3(_02813_),
    .B1(_02820_),
    .X(_00630_));
 sky130_fd_sc_hd__buf_2 _18616_ (.A(_05127_),
    .X(_02821_));
 sky130_fd_sc_hd__clkbuf_4 _18617_ (.A(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__xnor2_1 _18618_ (.A(_02822_),
    .B(\rbzero.wall_tracer.rayAddendY[2] ),
    .Y(_02823_));
 sky130_fd_sc_hd__a21oi_1 _18619_ (.A1(_02809_),
    .A2(_02813_),
    .B1(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__a311oi_1 _18620_ (.A1(_02809_),
    .A2(_02813_),
    .A3(_02823_),
    .B1(_02824_),
    .C1(_08136_),
    .Y(_02825_));
 sky130_fd_sc_hd__xor2_1 _18621_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(_05129_),
    .X(_02826_));
 sky130_fd_sc_hd__nor2_1 _18622_ (.A(_05132_),
    .B(\rbzero.debug_overlay.vplaneY[-8] ),
    .Y(_02827_));
 sky130_fd_sc_hd__and2b_1 _18623_ (.A_N(_02818_),
    .B(_02817_),
    .X(_02828_));
 sky130_fd_sc_hd__a21o_1 _18624_ (.A1(_02827_),
    .A2(_02816_),
    .B1(_02828_),
    .X(_02829_));
 sky130_fd_sc_hd__xnor2_1 _18625_ (.A(_02826_),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__xnor2_1 _18626_ (.A(_02814_),
    .B(_02830_),
    .Y(_02831_));
 sky130_fd_sc_hd__a21o_1 _18627_ (.A1(_02534_),
    .A2(_02831_),
    .B1(_09751_),
    .X(_02832_));
 sky130_fd_sc_hd__o22a_1 _18628_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(_02527_),
    .B1(_02825_),
    .B2(_02832_),
    .X(_00631_));
 sky130_fd_sc_hd__and2_1 _18629_ (.A(_05127_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_02833_));
 sky130_fd_sc_hd__nor2_1 _18630_ (.A(_05127_),
    .B(\rbzero.wall_tracer.rayAddendY[3] ),
    .Y(_02834_));
 sky130_fd_sc_hd__o21ai_1 _18631_ (.A1(\rbzero.wall_tracer.rayAddendY[2] ),
    .A2(\rbzero.wall_tracer.rayAddendY[1] ),
    .B1(_05127_),
    .Y(_02835_));
 sky130_fd_sc_hd__o21bai_1 _18632_ (.A1(_05127_),
    .A2(\rbzero.wall_tracer.rayAddendY[2] ),
    .B1_N(_02813_),
    .Y(_02836_));
 sky130_fd_sc_hd__o211ai_1 _18633_ (.A1(_02833_),
    .A2(_02834_),
    .B1(_02835_),
    .C1(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__a211o_1 _18634_ (.A1(_02835_),
    .A2(_02836_),
    .B1(_02833_),
    .C1(_02834_),
    .X(_02838_));
 sky130_fd_sc_hd__nand2_1 _18635_ (.A(_02826_),
    .B(_02829_),
    .Y(_02839_));
 sky130_fd_sc_hd__o21ai_1 _18636_ (.A1(_02828_),
    .A2(_02826_),
    .B1(_02814_),
    .Y(_02840_));
 sky130_fd_sc_hd__or2_1 _18637_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.debug_overlay.vplaneY[-5] ),
    .X(_02841_));
 sky130_fd_sc_hd__nand2_1 _18638_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(\rbzero.debug_overlay.vplaneY[-5] ),
    .Y(_02842_));
 sky130_fd_sc_hd__nand2_1 _18639_ (.A(_02841_),
    .B(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__or3_1 _18640_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(_05129_),
    .C(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__o21ai_1 _18641_ (.A1(\rbzero.debug_overlay.vplaneY[-2] ),
    .A2(_05129_),
    .B1(_02843_),
    .Y(_02845_));
 sky130_fd_sc_hd__nand2_1 _18642_ (.A(_02844_),
    .B(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__a21o_1 _18643_ (.A1(_02839_),
    .A2(_02840_),
    .B1(_02846_),
    .X(_02847_));
 sky130_fd_sc_hd__nand3_1 _18644_ (.A(_02839_),
    .B(_02846_),
    .C(_02840_),
    .Y(_02848_));
 sky130_fd_sc_hd__a32o_1 _18645_ (.A1(_08135_),
    .A2(_02847_),
    .A3(_02848_),
    .B1(_09751_),
    .B2(\rbzero.wall_tracer.rayAddendY[3] ),
    .X(_02849_));
 sky130_fd_sc_hd__a31o_1 _18646_ (.A1(_09753_),
    .A2(_02837_),
    .A3(_02838_),
    .B1(_02849_),
    .X(_00632_));
 sky130_fd_sc_hd__xor2_1 _18647_ (.A(_05127_),
    .B(\rbzero.wall_tracer.rayAddendY[4] ),
    .X(_02850_));
 sky130_fd_sc_hd__or2b_1 _18648_ (.A(_02833_),
    .B_N(_02838_),
    .X(_02851_));
 sky130_fd_sc_hd__xor2_1 _18649_ (.A(_02850_),
    .B(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__xnor2_1 _18650_ (.A(_02794_),
    .B(_05132_),
    .Y(_02853_));
 sky130_fd_sc_hd__a21o_1 _18651_ (.A1(_02844_),
    .A2(_02847_),
    .B1(_02853_),
    .X(_02854_));
 sky130_fd_sc_hd__nand3_1 _18652_ (.A(_02844_),
    .B(_02847_),
    .C(_02853_),
    .Y(_02855_));
 sky130_fd_sc_hd__a21oi_1 _18653_ (.A1(_02854_),
    .A2(_02855_),
    .B1(_02841_),
    .Y(_02856_));
 sky130_fd_sc_hd__a31o_1 _18654_ (.A1(_02841_),
    .A2(_02854_),
    .A3(_02855_),
    .B1(_04433_),
    .X(_02857_));
 sky130_fd_sc_hd__o22a_1 _18655_ (.A1(_08134_),
    .A2(_02852_),
    .B1(_02856_),
    .B2(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__mux2_1 _18656_ (.A0(\rbzero.wall_tracer.rayAddendY[4] ),
    .A1(_02858_),
    .S(_02525_),
    .X(_02859_));
 sky130_fd_sc_hd__clkbuf_1 _18657_ (.A(_02859_),
    .X(_00633_));
 sky130_fd_sc_hd__nand2_1 _18658_ (.A(_05127_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .Y(_02860_));
 sky130_fd_sc_hd__or2_1 _18659_ (.A(_05127_),
    .B(\rbzero.wall_tracer.rayAddendY[5] ),
    .X(_02861_));
 sky130_fd_sc_hd__nand2_1 _18660_ (.A(_02860_),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__or2b_1 _18661_ (.A(_02838_),
    .B_N(_02850_),
    .X(_02863_));
 sky130_fd_sc_hd__o21ai_1 _18662_ (.A1(\rbzero.wall_tracer.rayAddendY[4] ),
    .A2(\rbzero.wall_tracer.rayAddendY[3] ),
    .B1(_02821_),
    .Y(_02864_));
 sky130_fd_sc_hd__nand3_1 _18663_ (.A(_02862_),
    .B(_02863_),
    .C(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__a21o_1 _18664_ (.A1(_02863_),
    .A2(_02864_),
    .B1(_02862_),
    .X(_02866_));
 sky130_fd_sc_hd__a21o_1 _18665_ (.A1(_02847_),
    .A2(_02853_),
    .B1(_02841_),
    .X(_02867_));
 sky130_fd_sc_hd__nor2_1 _18666_ (.A(_02821_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .Y(_02868_));
 sky130_fd_sc_hd__and2_1 _18667_ (.A(_02821_),
    .B(\rbzero.debug_overlay.vplaneY[-3] ),
    .X(_02869_));
 sky130_fd_sc_hd__o22a_1 _18668_ (.A1(_02794_),
    .A2(_05132_),
    .B1(_02868_),
    .B2(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__nor4_1 _18669_ (.A(_02794_),
    .B(_05132_),
    .C(_02868_),
    .D(_02869_),
    .Y(_02871_));
 sky130_fd_sc_hd__or2_1 _18670_ (.A(_02870_),
    .B(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__a21oi_1 _18671_ (.A1(_02854_),
    .A2(_02867_),
    .B1(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__a31o_1 _18672_ (.A1(_02854_),
    .A2(_02872_),
    .A3(_02867_),
    .B1(_04434_),
    .X(_02874_));
 sky130_fd_sc_hd__a2bb2o_1 _18673_ (.A1_N(_02873_),
    .A2_N(_02874_),
    .B1(\rbzero.wall_tracer.rayAddendY[5] ),
    .B2(_09744_),
    .X(_02875_));
 sky130_fd_sc_hd__a31o_1 _18674_ (.A1(_09753_),
    .A2(_02865_),
    .A3(_02866_),
    .B1(_02875_),
    .X(_00634_));
 sky130_fd_sc_hd__xnor2_1 _18675_ (.A(_02821_),
    .B(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_02876_));
 sky130_fd_sc_hd__nand2_1 _18676_ (.A(_02860_),
    .B(_02866_),
    .Y(_02877_));
 sky130_fd_sc_hd__xnor2_1 _18677_ (.A(_02876_),
    .B(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__nor2_1 _18678_ (.A(_02821_),
    .B(\rbzero.debug_overlay.vplaneY[-2] ),
    .Y(_02879_));
 sky130_fd_sc_hd__and2_1 _18679_ (.A(_02821_),
    .B(\rbzero.debug_overlay.vplaneY[-2] ),
    .X(_02880_));
 sky130_fd_sc_hd__o21bai_1 _18680_ (.A1(_02879_),
    .A2(_02880_),
    .B1_N(_02868_),
    .Y(_02881_));
 sky130_fd_sc_hd__nand2_1 _18681_ (.A(\rbzero.debug_overlay.vplaneY[-2] ),
    .B(_02868_),
    .Y(_02882_));
 sky130_fd_sc_hd__nand2_1 _18682_ (.A(_02881_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__or2_1 _18683_ (.A(_02871_),
    .B(_02873_),
    .X(_02884_));
 sky130_fd_sc_hd__xnor2_1 _18684_ (.A(_02883_),
    .B(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__a22o_1 _18685_ (.A1(\rbzero.wall_tracer.rayAddendY[6] ),
    .A2(_09751_),
    .B1(_02885_),
    .B2(_08136_),
    .X(_02886_));
 sky130_fd_sc_hd__a21o_1 _18686_ (.A1(_09750_),
    .A2(_02878_),
    .B1(_02886_),
    .X(_00635_));
 sky130_fd_sc_hd__and2_1 _18687_ (.A(_02821_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_02887_));
 sky130_fd_sc_hd__nor2_1 _18688_ (.A(_02821_),
    .B(\rbzero.wall_tracer.rayAddendY[7] ),
    .Y(_02888_));
 sky130_fd_sc_hd__inv_2 _18689_ (.A(_02821_),
    .Y(_02889_));
 sky130_fd_sc_hd__inv_2 _18690_ (.A(\rbzero.wall_tracer.rayAddendY[6] ),
    .Y(_02890_));
 sky130_fd_sc_hd__or3_1 _18691_ (.A(_02862_),
    .B(_02863_),
    .C(_02876_),
    .X(_02891_));
 sky130_fd_sc_hd__o2111a_1 _18692_ (.A1(_02889_),
    .A2(_02890_),
    .B1(_02860_),
    .C1(_02864_),
    .D1(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__o21ai_1 _18693_ (.A1(_02887_),
    .A2(_02888_),
    .B1(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__or3_1 _18694_ (.A(_02887_),
    .B(_02888_),
    .C(_02892_),
    .X(_02894_));
 sky130_fd_sc_hd__nor2_1 _18695_ (.A(_02822_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .Y(_02895_));
 sky130_fd_sc_hd__and2_1 _18696_ (.A(_02822_),
    .B(\rbzero.debug_overlay.vplaneY[-1] ),
    .X(_02896_));
 sky130_fd_sc_hd__o21bai_1 _18697_ (.A1(_02895_),
    .A2(_02896_),
    .B1_N(_02879_),
    .Y(_02897_));
 sky130_fd_sc_hd__nand2_1 _18698_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_02879_),
    .Y(_02898_));
 sky130_fd_sc_hd__a21bo_1 _18699_ (.A1(_02881_),
    .A2(_02884_),
    .B1_N(_02882_),
    .X(_02899_));
 sky130_fd_sc_hd__nand3_1 _18700_ (.A(_02897_),
    .B(_02898_),
    .C(_02899_),
    .Y(_02900_));
 sky130_fd_sc_hd__a21o_1 _18701_ (.A1(_02897_),
    .A2(_02898_),
    .B1(_02899_),
    .X(_02901_));
 sky130_fd_sc_hd__a32o_1 _18702_ (.A1(_08135_),
    .A2(_02900_),
    .A3(_02901_),
    .B1(_09751_),
    .B2(\rbzero.wall_tracer.rayAddendY[7] ),
    .X(_02902_));
 sky130_fd_sc_hd__a31o_1 _18703_ (.A1(_09753_),
    .A2(_02893_),
    .A3(_02894_),
    .B1(_02902_),
    .X(_00636_));
 sky130_fd_sc_hd__xnor2_1 _18704_ (.A(_02822_),
    .B(\rbzero.wall_tracer.rayAddendY[8] ),
    .Y(_02903_));
 sky130_fd_sc_hd__and2b_1 _18705_ (.A_N(_02887_),
    .B(_02894_),
    .X(_02904_));
 sky130_fd_sc_hd__o21ai_1 _18706_ (.A1(_02903_),
    .A2(_02904_),
    .B1(_04434_),
    .Y(_02905_));
 sky130_fd_sc_hd__a21oi_1 _18707_ (.A1(_02903_),
    .A2(_02904_),
    .B1(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__inv_2 _18708_ (.A(_02794_),
    .Y(_02907_));
 sky130_fd_sc_hd__a21oi_1 _18709_ (.A1(_02794_),
    .A2(\rbzero.debug_overlay.vplaneY[-1] ),
    .B1(_02822_),
    .Y(_02908_));
 sky130_fd_sc_hd__a21oi_1 _18710_ (.A1(_02822_),
    .A2(_02794_),
    .B1(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__a21oi_1 _18711_ (.A1(_02907_),
    .A2(_02895_),
    .B1(_02909_),
    .Y(_02910_));
 sky130_fd_sc_hd__a21o_1 _18712_ (.A1(_02898_),
    .A2(_02900_),
    .B1(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__nand3_1 _18713_ (.A(_02898_),
    .B(_02900_),
    .C(_02910_),
    .Y(_02912_));
 sky130_fd_sc_hd__a31o_1 _18714_ (.A1(_08135_),
    .A2(_02911_),
    .A3(_02912_),
    .B1(_09745_),
    .X(_02913_));
 sky130_fd_sc_hd__o22a_1 _18715_ (.A1(\rbzero.wall_tracer.rayAddendY[8] ),
    .A2(_02527_),
    .B1(_02906_),
    .B2(_02913_),
    .X(_00637_));
 sky130_fd_sc_hd__or2_1 _18716_ (.A(_02822_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .X(_02914_));
 sky130_fd_sc_hd__nand2_1 _18717_ (.A(_02822_),
    .B(\rbzero.wall_tracer.rayAddendY[9] ),
    .Y(_02915_));
 sky130_fd_sc_hd__nand2_1 _18718_ (.A(_02914_),
    .B(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__nor2_1 _18719_ (.A(_02894_),
    .B(_02903_),
    .Y(_02917_));
 sky130_fd_sc_hd__a211o_1 _18720_ (.A1(_02822_),
    .A2(\rbzero.wall_tracer.rayAddendY[8] ),
    .B1(_02887_),
    .C1(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__xnor2_1 _18721_ (.A(_02916_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__a21oi_1 _18722_ (.A1(_02889_),
    .A2(_02907_),
    .B1(_02911_),
    .Y(_02920_));
 sky130_fd_sc_hd__a211o_1 _18723_ (.A1(_02908_),
    .A2(_02911_),
    .B1(_02920_),
    .C1(_04434_),
    .X(_02921_));
 sky130_fd_sc_hd__o221a_1 _18724_ (.A1(\rbzero.wall_tracer.rayAddendY[9] ),
    .A2(_02525_),
    .B1(_09760_),
    .B2(_02919_),
    .C1(_02921_),
    .X(_00638_));
 sky130_fd_sc_hd__a21bo_1 _18725_ (.A1(_02914_),
    .A2(_02918_),
    .B1_N(_02915_),
    .X(_02922_));
 sky130_fd_sc_hd__xnor2_1 _18726_ (.A(_02822_),
    .B(\rbzero.wall_tracer.rayAddendY[10] ),
    .Y(_02923_));
 sky130_fd_sc_hd__xnor2_1 _18727_ (.A(_02922_),
    .B(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__o21a_1 _18728_ (.A1(_02794_),
    .A2(_02911_),
    .B1(_08134_),
    .X(_02925_));
 sky130_fd_sc_hd__a22o_1 _18729_ (.A1(_04434_),
    .A2(_02924_),
    .B1(_02925_),
    .B2(_02889_),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_1 _18730_ (.A0(\rbzero.wall_tracer.rayAddendY[10] ),
    .A1(_02926_),
    .S(_02524_),
    .X(_02927_));
 sky130_fd_sc_hd__clkbuf_1 _18731_ (.A(_02927_),
    .X(_00639_));
 sky130_fd_sc_hd__and2b_1 _18732_ (.A_N(\rbzero.spi_registers.sclk_buffer[2] ),
    .B(\rbzero.spi_registers.sclk_buffer[1] ),
    .X(_02928_));
 sky130_fd_sc_hd__buf_2 _18733_ (.A(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__or2_2 _18734_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(\rbzero.spi_registers.spi_cmd[1] ),
    .X(_02930_));
 sky130_fd_sc_hd__a21o_1 _18735_ (.A1(\rbzero.spi_registers.spi_cmd[2] ),
    .A2(_02930_),
    .B1(\rbzero.spi_registers.spi_cmd[3] ),
    .X(_02931_));
 sky130_fd_sc_hd__nand2_1 _18736_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_02474_),
    .Y(_02932_));
 sky130_fd_sc_hd__and3b_1 _18737_ (.A_N(_02475_),
    .B(\rbzero.spi_registers.spi_cmd[3] ),
    .C(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__a31oi_2 _18738_ (.A1(_02474_),
    .A2(_02475_),
    .A3(_02476_),
    .B1(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__nand2_1 _18739_ (.A(_02931_),
    .B(_02934_),
    .Y(_02935_));
 sky130_fd_sc_hd__and2_1 _18740_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_02474_),
    .X(_02936_));
 sky130_fd_sc_hd__o21ai_1 _18741_ (.A1(_02475_),
    .A2(\rbzero.spi_registers.spi_cmd[3] ),
    .B1(\rbzero.spi_registers.spi_counter[2] ),
    .Y(_02937_));
 sky130_fd_sc_hd__o31a_1 _18742_ (.A1(\rbzero.spi_registers.spi_counter[2] ),
    .A2(_02475_),
    .A3(\rbzero.spi_registers.spi_cmd[3] ),
    .B1(\rbzero.spi_registers.spi_counter[1] ),
    .X(_02938_));
 sky130_fd_sc_hd__o211ai_1 _18743_ (.A1(_02936_),
    .A2(_02931_),
    .B1(_02937_),
    .C1(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__or4_1 _18744_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(\rbzero.spi_registers.spi_counter[1] ),
    .C(_02936_),
    .D(_02931_),
    .X(_02940_));
 sky130_fd_sc_hd__nand2_1 _18745_ (.A(_02939_),
    .B(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__nor3_1 _18746_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(\rbzero.spi_registers.spi_counter[0] ),
    .C(_02935_),
    .Y(_02942_));
 sky130_fd_sc_hd__a32o_1 _18747_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02935_),
    .A3(_02941_),
    .B1(_02942_),
    .B2(\rbzero.spi_registers.spi_counter[2] ),
    .X(_02943_));
 sky130_fd_sc_hd__or2_1 _18748_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02934_),
    .X(_02944_));
 sky130_fd_sc_hd__or2_1 _18749_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(\rbzero.spi_registers.spi_counter[5] ),
    .X(_02945_));
 sky130_fd_sc_hd__a21oi_1 _18750_ (.A1(\rbzero.spi_registers.spi_counter[4] ),
    .A2(_02934_),
    .B1(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hd__a31o_1 _18751_ (.A1(_02475_),
    .A2(_02932_),
    .A3(_02930_),
    .B1(\rbzero.spi_registers.spi_cmd[3] ),
    .X(_02947_));
 sky130_fd_sc_hd__or2b_1 _18752_ (.A(_02933_),
    .B_N(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__xnor2_1 _18753_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__and4_1 _18754_ (.A(_02943_),
    .B(_02944_),
    .C(_02946_),
    .D(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__nor2_2 _18755_ (.A(\rbzero.spi_registers.ss_buffer[1] ),
    .B(_04052_),
    .Y(_02951_));
 sky130_fd_sc_hd__a21bo_1 _18756_ (.A1(_02929_),
    .A2(_02950_),
    .B1_N(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__xnor2_1 _18757_ (.A(\rbzero.spi_registers.spi_counter[0] ),
    .B(_02929_),
    .Y(_02953_));
 sky130_fd_sc_hd__nor2_1 _18758_ (.A(_02952_),
    .B(_02953_),
    .Y(_00640_));
 sky130_fd_sc_hd__a21oi_1 _18759_ (.A1(\rbzero.spi_registers.spi_counter[0] ),
    .A2(_02929_),
    .B1(\rbzero.spi_registers.spi_counter[1] ),
    .Y(_02954_));
 sky130_fd_sc_hd__and3_1 _18760_ (.A(\rbzero.spi_registers.spi_counter[1] ),
    .B(\rbzero.spi_registers.spi_counter[0] ),
    .C(_02929_),
    .X(_02955_));
 sky130_fd_sc_hd__nor3_1 _18761_ (.A(_02952_),
    .B(_02954_),
    .C(_02955_),
    .Y(_00641_));
 sky130_fd_sc_hd__xnor2_1 _18762_ (.A(\rbzero.spi_registers.spi_counter[2] ),
    .B(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__nor2_1 _18763_ (.A(_02952_),
    .B(_02956_),
    .Y(_00642_));
 sky130_fd_sc_hd__and4_1 _18764_ (.A(\rbzero.spi_registers.spi_counter[3] ),
    .B(\rbzero.spi_registers.spi_counter[2] ),
    .C(\rbzero.spi_registers.spi_counter[1] ),
    .D(\rbzero.spi_registers.spi_counter[0] ),
    .X(_02957_));
 sky130_fd_sc_hd__a21oi_1 _18765_ (.A1(\rbzero.spi_registers.spi_counter[2] ),
    .A2(_02955_),
    .B1(\rbzero.spi_registers.spi_counter[3] ),
    .Y(_02958_));
 sky130_fd_sc_hd__a211oi_1 _18766_ (.A1(_02929_),
    .A2(_02957_),
    .B1(_02958_),
    .C1(_02952_),
    .Y(_00643_));
 sky130_fd_sc_hd__and3_1 _18767_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(_02929_),
    .C(_02957_),
    .X(_02959_));
 sky130_fd_sc_hd__a21oi_1 _18768_ (.A1(_02929_),
    .A2(_02957_),
    .B1(\rbzero.spi_registers.spi_counter[4] ),
    .Y(_02960_));
 sky130_fd_sc_hd__nor3_1 _18769_ (.A(_02952_),
    .B(_02959_),
    .C(_02960_),
    .Y(_00644_));
 sky130_fd_sc_hd__and2_1 _18770_ (.A(\rbzero.spi_registers.spi_counter[5] ),
    .B(_02959_),
    .X(_02961_));
 sky130_fd_sc_hd__o21ai_1 _18771_ (.A1(\rbzero.spi_registers.spi_counter[5] ),
    .A2(_02959_),
    .B1(_02951_),
    .Y(_02962_));
 sky130_fd_sc_hd__nor2_1 _18772_ (.A(_02961_),
    .B(_02962_),
    .Y(_00645_));
 sky130_fd_sc_hd__or2_1 _18773_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(_02961_),
    .X(_02963_));
 sky130_fd_sc_hd__nand2_1 _18774_ (.A(\rbzero.spi_registers.spi_counter[6] ),
    .B(_02961_),
    .Y(_02964_));
 sky130_fd_sc_hd__and3_1 _18775_ (.A(_02951_),
    .B(_02963_),
    .C(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__clkbuf_1 _18776_ (.A(_02965_),
    .X(_00646_));
 sky130_fd_sc_hd__nand2_1 _18777_ (.A(\rbzero.pov.spi_done ),
    .B(_08116_),
    .Y(_02966_));
 sky130_fd_sc_hd__buf_4 _18778_ (.A(_02966_),
    .X(_02967_));
 sky130_fd_sc_hd__buf_4 _18779_ (.A(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__mux2_1 _18780_ (.A0(\rbzero.pov.spi_buffer[0] ),
    .A1(\rbzero.pov.ready_buffer[0] ),
    .S(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__clkbuf_1 _18781_ (.A(_02969_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _18782_ (.A0(\rbzero.pov.spi_buffer[1] ),
    .A1(\rbzero.pov.ready_buffer[1] ),
    .S(_02968_),
    .X(_02970_));
 sky130_fd_sc_hd__clkbuf_1 _18783_ (.A(_02970_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _18784_ (.A0(\rbzero.pov.spi_buffer[2] ),
    .A1(\rbzero.pov.ready_buffer[2] ),
    .S(_02968_),
    .X(_02971_));
 sky130_fd_sc_hd__clkbuf_1 _18785_ (.A(_02971_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _18786_ (.A0(\rbzero.pov.spi_buffer[3] ),
    .A1(\rbzero.pov.ready_buffer[3] ),
    .S(_02968_),
    .X(_02972_));
 sky130_fd_sc_hd__clkbuf_1 _18787_ (.A(_02972_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _18788_ (.A0(\rbzero.pov.spi_buffer[4] ),
    .A1(\rbzero.pov.ready_buffer[4] ),
    .S(_02968_),
    .X(_02973_));
 sky130_fd_sc_hd__clkbuf_1 _18789_ (.A(_02973_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _18790_ (.A0(\rbzero.pov.spi_buffer[5] ),
    .A1(\rbzero.pov.ready_buffer[5] ),
    .S(_02968_),
    .X(_02974_));
 sky130_fd_sc_hd__clkbuf_1 _18791_ (.A(_02974_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _18792_ (.A0(\rbzero.pov.spi_buffer[6] ),
    .A1(\rbzero.pov.ready_buffer[6] ),
    .S(_02968_),
    .X(_02975_));
 sky130_fd_sc_hd__clkbuf_1 _18793_ (.A(_02975_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _18794_ (.A0(\rbzero.pov.spi_buffer[7] ),
    .A1(\rbzero.pov.ready_buffer[7] ),
    .S(_02968_),
    .X(_02976_));
 sky130_fd_sc_hd__clkbuf_1 _18795_ (.A(_02976_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _18796_ (.A0(\rbzero.pov.spi_buffer[8] ),
    .A1(\rbzero.pov.ready_buffer[8] ),
    .S(_02968_),
    .X(_02977_));
 sky130_fd_sc_hd__clkbuf_1 _18797_ (.A(_02977_),
    .X(_00655_));
 sky130_fd_sc_hd__clkbuf_4 _18798_ (.A(_02967_),
    .X(_02978_));
 sky130_fd_sc_hd__mux2_1 _18799_ (.A0(\rbzero.pov.spi_buffer[9] ),
    .A1(\rbzero.pov.ready_buffer[9] ),
    .S(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__clkbuf_1 _18800_ (.A(_02979_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _18801_ (.A0(\rbzero.pov.spi_buffer[10] ),
    .A1(\rbzero.pov.ready_buffer[10] ),
    .S(_02978_),
    .X(_02980_));
 sky130_fd_sc_hd__clkbuf_1 _18802_ (.A(_02980_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _18803_ (.A0(\rbzero.pov.spi_buffer[11] ),
    .A1(\rbzero.pov.ready_buffer[11] ),
    .S(_02978_),
    .X(_02981_));
 sky130_fd_sc_hd__clkbuf_1 _18804_ (.A(_02981_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _18805_ (.A0(\rbzero.pov.spi_buffer[12] ),
    .A1(\rbzero.pov.ready_buffer[12] ),
    .S(_02978_),
    .X(_02982_));
 sky130_fd_sc_hd__clkbuf_1 _18806_ (.A(_02982_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _18807_ (.A0(\rbzero.pov.spi_buffer[13] ),
    .A1(\rbzero.pov.ready_buffer[13] ),
    .S(_02978_),
    .X(_02983_));
 sky130_fd_sc_hd__clkbuf_1 _18808_ (.A(_02983_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _18809_ (.A0(\rbzero.pov.spi_buffer[14] ),
    .A1(\rbzero.pov.ready_buffer[14] ),
    .S(_02978_),
    .X(_02984_));
 sky130_fd_sc_hd__clkbuf_1 _18810_ (.A(_02984_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _18811_ (.A0(\rbzero.pov.spi_buffer[15] ),
    .A1(\rbzero.pov.ready_buffer[15] ),
    .S(_02978_),
    .X(_02985_));
 sky130_fd_sc_hd__clkbuf_1 _18812_ (.A(_02985_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _18813_ (.A0(\rbzero.pov.spi_buffer[16] ),
    .A1(\rbzero.pov.ready_buffer[16] ),
    .S(_02978_),
    .X(_02986_));
 sky130_fd_sc_hd__clkbuf_1 _18814_ (.A(_02986_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _18815_ (.A0(\rbzero.pov.spi_buffer[17] ),
    .A1(\rbzero.pov.ready_buffer[17] ),
    .S(_02978_),
    .X(_02987_));
 sky130_fd_sc_hd__clkbuf_1 _18816_ (.A(_02987_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _18817_ (.A0(\rbzero.pov.spi_buffer[18] ),
    .A1(\rbzero.pov.ready_buffer[18] ),
    .S(_02978_),
    .X(_02988_));
 sky130_fd_sc_hd__clkbuf_1 _18818_ (.A(_02988_),
    .X(_00665_));
 sky130_fd_sc_hd__clkbuf_4 _18819_ (.A(_02967_),
    .X(_02989_));
 sky130_fd_sc_hd__mux2_1 _18820_ (.A0(\rbzero.pov.spi_buffer[19] ),
    .A1(\rbzero.pov.ready_buffer[19] ),
    .S(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__clkbuf_1 _18821_ (.A(_02990_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _18822_ (.A0(\rbzero.pov.spi_buffer[20] ),
    .A1(\rbzero.pov.ready_buffer[20] ),
    .S(_02989_),
    .X(_02991_));
 sky130_fd_sc_hd__clkbuf_1 _18823_ (.A(_02991_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _18824_ (.A0(\rbzero.pov.spi_buffer[21] ),
    .A1(\rbzero.pov.ready_buffer[21] ),
    .S(_02989_),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_1 _18825_ (.A(_02992_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _18826_ (.A0(\rbzero.pov.spi_buffer[22] ),
    .A1(\rbzero.pov.ready_buffer[22] ),
    .S(_02989_),
    .X(_02993_));
 sky130_fd_sc_hd__clkbuf_1 _18827_ (.A(_02993_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _18828_ (.A0(\rbzero.pov.spi_buffer[23] ),
    .A1(\rbzero.pov.ready_buffer[23] ),
    .S(_02989_),
    .X(_02994_));
 sky130_fd_sc_hd__clkbuf_1 _18829_ (.A(_02994_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _18830_ (.A0(\rbzero.pov.spi_buffer[24] ),
    .A1(\rbzero.pov.ready_buffer[24] ),
    .S(_02989_),
    .X(_02995_));
 sky130_fd_sc_hd__clkbuf_1 _18831_ (.A(_02995_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _18832_ (.A0(\rbzero.pov.spi_buffer[25] ),
    .A1(\rbzero.pov.ready_buffer[25] ),
    .S(_02989_),
    .X(_02996_));
 sky130_fd_sc_hd__clkbuf_1 _18833_ (.A(_02996_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _18834_ (.A0(\rbzero.pov.spi_buffer[26] ),
    .A1(\rbzero.pov.ready_buffer[26] ),
    .S(_02989_),
    .X(_02997_));
 sky130_fd_sc_hd__clkbuf_1 _18835_ (.A(_02997_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _18836_ (.A0(\rbzero.pov.spi_buffer[27] ),
    .A1(\rbzero.pov.ready_buffer[27] ),
    .S(_02989_),
    .X(_02998_));
 sky130_fd_sc_hd__clkbuf_1 _18837_ (.A(_02998_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _18838_ (.A0(\rbzero.pov.spi_buffer[28] ),
    .A1(\rbzero.pov.ready_buffer[28] ),
    .S(_02989_),
    .X(_02999_));
 sky130_fd_sc_hd__clkbuf_1 _18839_ (.A(_02999_),
    .X(_00675_));
 sky130_fd_sc_hd__clkbuf_4 _18840_ (.A(_02967_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_1 _18841_ (.A0(\rbzero.pov.spi_buffer[29] ),
    .A1(\rbzero.pov.ready_buffer[29] ),
    .S(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__clkbuf_1 _18842_ (.A(_03001_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _18843_ (.A0(\rbzero.pov.spi_buffer[30] ),
    .A1(\rbzero.pov.ready_buffer[30] ),
    .S(_03000_),
    .X(_03002_));
 sky130_fd_sc_hd__clkbuf_1 _18844_ (.A(_03002_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _18845_ (.A0(\rbzero.pov.spi_buffer[31] ),
    .A1(\rbzero.pov.ready_buffer[31] ),
    .S(_03000_),
    .X(_03003_));
 sky130_fd_sc_hd__clkbuf_1 _18846_ (.A(_03003_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _18847_ (.A0(\rbzero.pov.spi_buffer[32] ),
    .A1(\rbzero.pov.ready_buffer[32] ),
    .S(_03000_),
    .X(_03004_));
 sky130_fd_sc_hd__clkbuf_1 _18848_ (.A(_03004_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _18849_ (.A0(\rbzero.pov.spi_buffer[33] ),
    .A1(\rbzero.pov.ready_buffer[33] ),
    .S(_03000_),
    .X(_03005_));
 sky130_fd_sc_hd__clkbuf_1 _18850_ (.A(_03005_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _18851_ (.A0(\rbzero.pov.spi_buffer[34] ),
    .A1(\rbzero.pov.ready_buffer[34] ),
    .S(_03000_),
    .X(_03006_));
 sky130_fd_sc_hd__clkbuf_1 _18852_ (.A(_03006_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _18853_ (.A0(\rbzero.pov.spi_buffer[35] ),
    .A1(\rbzero.pov.ready_buffer[35] ),
    .S(_03000_),
    .X(_03007_));
 sky130_fd_sc_hd__clkbuf_1 _18854_ (.A(_03007_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _18855_ (.A0(\rbzero.pov.spi_buffer[36] ),
    .A1(\rbzero.pov.ready_buffer[36] ),
    .S(_03000_),
    .X(_03008_));
 sky130_fd_sc_hd__clkbuf_1 _18856_ (.A(_03008_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _18857_ (.A0(\rbzero.pov.spi_buffer[37] ),
    .A1(\rbzero.pov.ready_buffer[37] ),
    .S(_03000_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_1 _18858_ (.A(_03009_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _18859_ (.A0(\rbzero.pov.spi_buffer[38] ),
    .A1(\rbzero.pov.ready_buffer[38] ),
    .S(_03000_),
    .X(_03010_));
 sky130_fd_sc_hd__clkbuf_1 _18860_ (.A(_03010_),
    .X(_00685_));
 sky130_fd_sc_hd__buf_4 _18861_ (.A(_02967_),
    .X(_03011_));
 sky130_fd_sc_hd__mux2_1 _18862_ (.A0(\rbzero.pov.spi_buffer[39] ),
    .A1(\rbzero.pov.ready_buffer[39] ),
    .S(_03011_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_1 _18863_ (.A(_03012_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _18864_ (.A0(\rbzero.pov.spi_buffer[40] ),
    .A1(\rbzero.pov.ready_buffer[40] ),
    .S(_03011_),
    .X(_03013_));
 sky130_fd_sc_hd__clkbuf_1 _18865_ (.A(_03013_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _18866_ (.A0(\rbzero.pov.spi_buffer[41] ),
    .A1(\rbzero.pov.ready_buffer[41] ),
    .S(_03011_),
    .X(_03014_));
 sky130_fd_sc_hd__clkbuf_1 _18867_ (.A(_03014_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _18868_ (.A0(\rbzero.pov.spi_buffer[42] ),
    .A1(\rbzero.pov.ready_buffer[42] ),
    .S(_03011_),
    .X(_03015_));
 sky130_fd_sc_hd__clkbuf_1 _18869_ (.A(_03015_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _18870_ (.A0(\rbzero.pov.spi_buffer[43] ),
    .A1(\rbzero.pov.ready_buffer[43] ),
    .S(_03011_),
    .X(_03016_));
 sky130_fd_sc_hd__clkbuf_1 _18871_ (.A(_03016_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _18872_ (.A0(\rbzero.pov.spi_buffer[44] ),
    .A1(\rbzero.pov.ready_buffer[44] ),
    .S(_03011_),
    .X(_03017_));
 sky130_fd_sc_hd__clkbuf_1 _18873_ (.A(_03017_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _18874_ (.A0(\rbzero.pov.spi_buffer[45] ),
    .A1(\rbzero.pov.ready_buffer[45] ),
    .S(_03011_),
    .X(_03018_));
 sky130_fd_sc_hd__clkbuf_1 _18875_ (.A(_03018_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _18876_ (.A0(\rbzero.pov.spi_buffer[46] ),
    .A1(\rbzero.pov.ready_buffer[46] ),
    .S(_03011_),
    .X(_03019_));
 sky130_fd_sc_hd__clkbuf_1 _18877_ (.A(_03019_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _18878_ (.A0(\rbzero.pov.spi_buffer[47] ),
    .A1(\rbzero.pov.ready_buffer[47] ),
    .S(_03011_),
    .X(_03020_));
 sky130_fd_sc_hd__clkbuf_1 _18879_ (.A(_03020_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _18880_ (.A0(\rbzero.pov.spi_buffer[48] ),
    .A1(\rbzero.pov.ready_buffer[48] ),
    .S(_03011_),
    .X(_03021_));
 sky130_fd_sc_hd__clkbuf_1 _18881_ (.A(_03021_),
    .X(_00695_));
 sky130_fd_sc_hd__buf_4 _18882_ (.A(_02966_),
    .X(_03022_));
 sky130_fd_sc_hd__mux2_1 _18883_ (.A0(\rbzero.pov.spi_buffer[49] ),
    .A1(\rbzero.pov.ready_buffer[49] ),
    .S(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__clkbuf_1 _18884_ (.A(_03023_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _18885_ (.A0(\rbzero.pov.spi_buffer[50] ),
    .A1(\rbzero.pov.ready_buffer[50] ),
    .S(_03022_),
    .X(_03024_));
 sky130_fd_sc_hd__clkbuf_1 _18886_ (.A(_03024_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _18887_ (.A0(\rbzero.pov.spi_buffer[51] ),
    .A1(\rbzero.pov.ready_buffer[51] ),
    .S(_03022_),
    .X(_03025_));
 sky130_fd_sc_hd__clkbuf_1 _18888_ (.A(_03025_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _18889_ (.A0(\rbzero.pov.spi_buffer[52] ),
    .A1(\rbzero.pov.ready_buffer[52] ),
    .S(_03022_),
    .X(_03026_));
 sky130_fd_sc_hd__clkbuf_1 _18890_ (.A(_03026_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _18891_ (.A0(\rbzero.pov.spi_buffer[53] ),
    .A1(\rbzero.pov.ready_buffer[53] ),
    .S(_03022_),
    .X(_03027_));
 sky130_fd_sc_hd__clkbuf_1 _18892_ (.A(_03027_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _18893_ (.A0(\rbzero.pov.spi_buffer[54] ),
    .A1(\rbzero.pov.ready_buffer[54] ),
    .S(_03022_),
    .X(_03028_));
 sky130_fd_sc_hd__clkbuf_1 _18894_ (.A(_03028_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _18895_ (.A0(\rbzero.pov.spi_buffer[55] ),
    .A1(\rbzero.pov.ready_buffer[55] ),
    .S(_03022_),
    .X(_03029_));
 sky130_fd_sc_hd__clkbuf_1 _18896_ (.A(_03029_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _18897_ (.A0(\rbzero.pov.spi_buffer[56] ),
    .A1(\rbzero.pov.ready_buffer[56] ),
    .S(_03022_),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_1 _18898_ (.A(_03030_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _18899_ (.A0(\rbzero.pov.spi_buffer[57] ),
    .A1(\rbzero.pov.ready_buffer[57] ),
    .S(_03022_),
    .X(_03031_));
 sky130_fd_sc_hd__clkbuf_1 _18900_ (.A(_03031_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _18901_ (.A0(\rbzero.pov.spi_buffer[58] ),
    .A1(\rbzero.pov.ready_buffer[58] ),
    .S(_03022_),
    .X(_03032_));
 sky130_fd_sc_hd__clkbuf_1 _18902_ (.A(_03032_),
    .X(_00705_));
 sky130_fd_sc_hd__buf_4 _18903_ (.A(_02966_),
    .X(_03033_));
 sky130_fd_sc_hd__mux2_1 _18904_ (.A0(\rbzero.pov.spi_buffer[59] ),
    .A1(\rbzero.pov.ready_buffer[59] ),
    .S(_03033_),
    .X(_03034_));
 sky130_fd_sc_hd__clkbuf_1 _18905_ (.A(_03034_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _18906_ (.A0(\rbzero.pov.spi_buffer[60] ),
    .A1(\rbzero.pov.ready_buffer[60] ),
    .S(_03033_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_1 _18907_ (.A(_03035_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _18908_ (.A0(\rbzero.pov.spi_buffer[61] ),
    .A1(\rbzero.pov.ready_buffer[61] ),
    .S(_03033_),
    .X(_03036_));
 sky130_fd_sc_hd__clkbuf_1 _18909_ (.A(_03036_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _18910_ (.A0(\rbzero.pov.spi_buffer[62] ),
    .A1(\rbzero.pov.ready_buffer[62] ),
    .S(_03033_),
    .X(_03037_));
 sky130_fd_sc_hd__clkbuf_1 _18911_ (.A(_03037_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _18912_ (.A0(\rbzero.pov.spi_buffer[63] ),
    .A1(\rbzero.pov.ready_buffer[63] ),
    .S(_03033_),
    .X(_03038_));
 sky130_fd_sc_hd__clkbuf_1 _18913_ (.A(_03038_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _18914_ (.A0(\rbzero.pov.spi_buffer[64] ),
    .A1(\rbzero.pov.ready_buffer[64] ),
    .S(_03033_),
    .X(_03039_));
 sky130_fd_sc_hd__clkbuf_1 _18915_ (.A(_03039_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _18916_ (.A0(\rbzero.pov.spi_buffer[65] ),
    .A1(\rbzero.pov.ready_buffer[65] ),
    .S(_03033_),
    .X(_03040_));
 sky130_fd_sc_hd__clkbuf_1 _18917_ (.A(_03040_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _18918_ (.A0(\rbzero.pov.spi_buffer[66] ),
    .A1(\rbzero.pov.ready_buffer[66] ),
    .S(_03033_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_1 _18919_ (.A(_03041_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _18920_ (.A0(\rbzero.pov.spi_buffer[67] ),
    .A1(\rbzero.pov.ready_buffer[67] ),
    .S(_03033_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _18921_ (.A(_03042_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _18922_ (.A0(\rbzero.pov.spi_buffer[68] ),
    .A1(\rbzero.pov.ready_buffer[68] ),
    .S(_03033_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _18923_ (.A(_03043_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _18924_ (.A0(\rbzero.pov.spi_buffer[69] ),
    .A1(\rbzero.pov.ready_buffer[69] ),
    .S(_02967_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_1 _18925_ (.A(_03044_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _18926_ (.A0(\rbzero.pov.spi_buffer[70] ),
    .A1(\rbzero.pov.ready_buffer[70] ),
    .S(_02967_),
    .X(_03045_));
 sky130_fd_sc_hd__clkbuf_1 _18927_ (.A(_03045_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _18928_ (.A0(\rbzero.pov.spi_buffer[71] ),
    .A1(\rbzero.pov.ready_buffer[71] ),
    .S(_02967_),
    .X(_03046_));
 sky130_fd_sc_hd__clkbuf_1 _18929_ (.A(_03046_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _18930_ (.A0(\rbzero.pov.spi_buffer[72] ),
    .A1(\rbzero.pov.ready_buffer[72] ),
    .S(_02967_),
    .X(_03047_));
 sky130_fd_sc_hd__clkbuf_1 _18931_ (.A(_03047_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _18932_ (.A0(\rbzero.pov.spi_buffer[73] ),
    .A1(\rbzero.pov.ready_buffer[73] ),
    .S(_02967_),
    .X(_03048_));
 sky130_fd_sc_hd__clkbuf_1 _18933_ (.A(_03048_),
    .X(_00720_));
 sky130_fd_sc_hd__nor4_1 _18934_ (.A(\rbzero.spi_registers.spi_counter[4] ),
    .B(\rbzero.spi_registers.spi_counter[3] ),
    .C(\rbzero.spi_registers.spi_counter[2] ),
    .D(_02945_),
    .Y(_03049_));
 sky130_fd_sc_hd__and3b_1 _18935_ (.A_N(_03049_),
    .B(_02929_),
    .C(_02951_),
    .X(_03050_));
 sky130_fd_sc_hd__clkbuf_4 _18936_ (.A(_03050_),
    .X(_03051_));
 sky130_fd_sc_hd__buf_4 _18937_ (.A(_03051_),
    .X(_03052_));
 sky130_fd_sc_hd__mux2_1 _18938_ (.A0(_02473_),
    .A1(\rbzero.spi_registers.mosi ),
    .S(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__clkbuf_1 _18939_ (.A(_03053_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _18940_ (.A0(_02481_),
    .A1(_02473_),
    .S(_03052_),
    .X(_03054_));
 sky130_fd_sc_hd__clkbuf_1 _18941_ (.A(_03054_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _18942_ (.A0(_02483_),
    .A1(_02481_),
    .S(_03052_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_1 _18943_ (.A(_03055_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _18944_ (.A0(_02485_),
    .A1(_02483_),
    .S(_03052_),
    .X(_03056_));
 sky130_fd_sc_hd__clkbuf_1 _18945_ (.A(_03056_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _18946_ (.A0(_02487_),
    .A1(_02485_),
    .S(_03052_),
    .X(_03057_));
 sky130_fd_sc_hd__clkbuf_1 _18947_ (.A(_03057_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _18948_ (.A0(_02489_),
    .A1(_02487_),
    .S(_03052_),
    .X(_03058_));
 sky130_fd_sc_hd__clkbuf_1 _18949_ (.A(_03058_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _18950_ (.A0(\rbzero.spi_registers.spi_buffer[6] ),
    .A1(_02489_),
    .S(_03052_),
    .X(_03059_));
 sky130_fd_sc_hd__clkbuf_1 _18951_ (.A(_03059_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _18952_ (.A0(\rbzero.spi_registers.spi_buffer[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03052_),
    .X(_03060_));
 sky130_fd_sc_hd__clkbuf_1 _18953_ (.A(_03060_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _18954_ (.A0(\rbzero.spi_registers.spi_buffer[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03052_),
    .X(_03061_));
 sky130_fd_sc_hd__clkbuf_1 _18955_ (.A(_03061_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _18956_ (.A0(\rbzero.spi_registers.spi_buffer[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03052_),
    .X(_03062_));
 sky130_fd_sc_hd__clkbuf_1 _18957_ (.A(_03062_),
    .X(_00730_));
 sky130_fd_sc_hd__buf_4 _18958_ (.A(_03051_),
    .X(_03063_));
 sky130_fd_sc_hd__mux2_1 _18959_ (.A0(\rbzero.spi_registers.spi_buffer[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__clkbuf_1 _18960_ (.A(_03064_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _18961_ (.A0(\rbzero.spi_registers.spi_buffer[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03063_),
    .X(_03065_));
 sky130_fd_sc_hd__clkbuf_1 _18962_ (.A(_03065_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _18963_ (.A0(\rbzero.spi_registers.spi_buffer[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03063_),
    .X(_03066_));
 sky130_fd_sc_hd__clkbuf_1 _18964_ (.A(_03066_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _18965_ (.A0(\rbzero.spi_registers.spi_buffer[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03063_),
    .X(_03067_));
 sky130_fd_sc_hd__clkbuf_1 _18966_ (.A(_03067_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _18967_ (.A0(\rbzero.spi_registers.spi_buffer[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03063_),
    .X(_03068_));
 sky130_fd_sc_hd__clkbuf_1 _18968_ (.A(_03068_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _18969_ (.A0(\rbzero.spi_registers.spi_buffer[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03063_),
    .X(_03069_));
 sky130_fd_sc_hd__clkbuf_1 _18970_ (.A(_03069_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _18971_ (.A0(\rbzero.spi_registers.spi_buffer[16] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03063_),
    .X(_03070_));
 sky130_fd_sc_hd__clkbuf_1 _18972_ (.A(_03070_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _18973_ (.A0(\rbzero.spi_registers.spi_buffer[17] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03063_),
    .X(_03071_));
 sky130_fd_sc_hd__clkbuf_1 _18974_ (.A(_03071_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _18975_ (.A0(\rbzero.spi_registers.spi_buffer[18] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03063_),
    .X(_03072_));
 sky130_fd_sc_hd__clkbuf_1 _18976_ (.A(_03072_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _18977_ (.A0(\rbzero.spi_registers.spi_buffer[19] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03063_),
    .X(_03073_));
 sky130_fd_sc_hd__clkbuf_1 _18978_ (.A(_03073_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _18979_ (.A0(\rbzero.spi_registers.spi_buffer[20] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03051_),
    .X(_03074_));
 sky130_fd_sc_hd__clkbuf_1 _18980_ (.A(_03074_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _18981_ (.A0(\rbzero.spi_registers.spi_buffer[21] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03051_),
    .X(_03075_));
 sky130_fd_sc_hd__clkbuf_1 _18982_ (.A(_03075_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _18983_ (.A0(\rbzero.spi_registers.spi_buffer[22] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03051_),
    .X(_03076_));
 sky130_fd_sc_hd__clkbuf_1 _18984_ (.A(_03076_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _18985_ (.A0(\rbzero.spi_registers.spi_buffer[23] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03051_),
    .X(_03077_));
 sky130_fd_sc_hd__clkbuf_1 _18986_ (.A(_03077_),
    .X(_00744_));
 sky130_fd_sc_hd__and3_1 _18987_ (.A(_02951_),
    .B(_02929_),
    .C(_03049_),
    .X(_03078_));
 sky130_fd_sc_hd__mux2_1 _18988_ (.A0(\rbzero.spi_registers.spi_cmd[0] ),
    .A1(\rbzero.spi_registers.mosi ),
    .S(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__clkbuf_1 _18989_ (.A(_03079_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _18990_ (.A0(_02474_),
    .A1(\rbzero.spi_registers.spi_cmd[0] ),
    .S(_03078_),
    .X(_03080_));
 sky130_fd_sc_hd__clkbuf_1 _18991_ (.A(_03080_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _18992_ (.A0(_02475_),
    .A1(_02474_),
    .S(_03078_),
    .X(_03081_));
 sky130_fd_sc_hd__clkbuf_1 _18993_ (.A(_03081_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _18994_ (.A0(\rbzero.spi_registers.spi_cmd[3] ),
    .A1(_02475_),
    .S(_03078_),
    .X(_03082_));
 sky130_fd_sc_hd__clkbuf_1 _18995_ (.A(_03082_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _18996_ (.A0(net44),
    .A1(\rbzero.spi_registers.mosi_buffer[0] ),
    .S(_09734_),
    .X(_03083_));
 sky130_fd_sc_hd__clkbuf_1 _18997_ (.A(_03083_),
    .X(_00749_));
 sky130_fd_sc_hd__clkbuf_4 _18998_ (.A(_08116_),
    .X(_03084_));
 sky130_fd_sc_hd__mux2_1 _18999_ (.A0(\rbzero.spi_registers.mosi ),
    .A1(\rbzero.spi_registers.mosi_buffer[0] ),
    .S(_03084_),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_1 _19000_ (.A(_03085_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _19001_ (.A0(net43),
    .A1(\rbzero.spi_registers.ss_buffer[0] ),
    .S(_09734_),
    .X(_03086_));
 sky130_fd_sc_hd__clkbuf_1 _19002_ (.A(_03086_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _19003_ (.A0(\rbzero.spi_registers.ss_buffer[1] ),
    .A1(\rbzero.spi_registers.ss_buffer[0] ),
    .S(_03084_),
    .X(_03087_));
 sky130_fd_sc_hd__clkbuf_1 _19004_ (.A(_03087_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _19005_ (.A0(net46),
    .A1(\rbzero.spi_registers.sclk_buffer[0] ),
    .S(_09734_),
    .X(_03088_));
 sky130_fd_sc_hd__clkbuf_1 _19006_ (.A(_03088_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _19007_ (.A0(\rbzero.spi_registers.sclk_buffer[1] ),
    .A1(\rbzero.spi_registers.sclk_buffer[0] ),
    .S(_03084_),
    .X(_03089_));
 sky130_fd_sc_hd__clkbuf_1 _19008_ (.A(_03089_),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _19009_ (.A0(\rbzero.spi_registers.sclk_buffer[2] ),
    .A1(\rbzero.spi_registers.sclk_buffer[1] ),
    .S(_03084_),
    .X(_03090_));
 sky130_fd_sc_hd__clkbuf_1 _19010_ (.A(_03090_),
    .X(_00755_));
 sky130_fd_sc_hd__and4b_2 _19011_ (.A_N(_05653_),
    .B(_05652_),
    .C(_04642_),
    .D(_05645_),
    .X(_03091_));
 sky130_fd_sc_hd__and3_1 _19012_ (.A(_04687_),
    .B(_05651_),
    .C(\gpout0.vpos[0] ),
    .X(_03092_));
 sky130_fd_sc_hd__and3_1 _19013_ (.A(_05644_),
    .B(_09747_),
    .C(_03092_),
    .X(_03093_));
 sky130_fd_sc_hd__and3_1 _19014_ (.A(_05270_),
    .B(_03091_),
    .C(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__buf_6 _19015_ (.A(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__buf_6 _19016_ (.A(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__buf_4 _19017_ (.A(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__nand2_4 _19018_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__and3_1 _19019_ (.A(_05644_),
    .B(_09728_),
    .C(_03092_),
    .X(_03099_));
 sky130_fd_sc_hd__and3_4 _19020_ (.A(_05270_),
    .B(_03091_),
    .C(_03099_),
    .X(_03100_));
 sky130_fd_sc_hd__and2_2 _19021_ (.A(\rbzero.spi_registers.got_new_other ),
    .B(_03100_),
    .X(_03101_));
 sky130_fd_sc_hd__or2_1 _19022_ (.A(\rbzero.map_overlay.i_otherx[0] ),
    .B(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__clkbuf_4 _19023_ (.A(_03084_),
    .X(_03103_));
 sky130_fd_sc_hd__o211a_1 _19024_ (.A1(\rbzero.spi_registers.new_other[6] ),
    .A2(_03098_),
    .B1(_03102_),
    .C1(_03103_),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _19025_ (.A(\rbzero.map_overlay.i_otherx[1] ),
    .B(_03101_),
    .X(_03104_));
 sky130_fd_sc_hd__o211a_1 _19026_ (.A1(\rbzero.spi_registers.new_other[7] ),
    .A2(_03098_),
    .B1(_03104_),
    .C1(_03103_),
    .X(_00757_));
 sky130_fd_sc_hd__or2_1 _19027_ (.A(\rbzero.map_overlay.i_otherx[2] ),
    .B(_03101_),
    .X(_03105_));
 sky130_fd_sc_hd__o211a_1 _19028_ (.A1(\rbzero.spi_registers.new_other[8] ),
    .A2(_03098_),
    .B1(_03105_),
    .C1(_03103_),
    .X(_00758_));
 sky130_fd_sc_hd__or2_1 _19029_ (.A(\rbzero.map_overlay.i_otherx[3] ),
    .B(_03101_),
    .X(_03106_));
 sky130_fd_sc_hd__o211a_1 _19030_ (.A1(\rbzero.spi_registers.new_other[9] ),
    .A2(_03098_),
    .B1(_03106_),
    .C1(_03103_),
    .X(_00759_));
 sky130_fd_sc_hd__or2_1 _19031_ (.A(\rbzero.map_overlay.i_otherx[4] ),
    .B(_03101_),
    .X(_03107_));
 sky130_fd_sc_hd__o211a_1 _19032_ (.A1(\rbzero.spi_registers.new_other[10] ),
    .A2(_03098_),
    .B1(_03107_),
    .C1(_03103_),
    .X(_00760_));
 sky130_fd_sc_hd__or2_1 _19033_ (.A(\rbzero.map_overlay.i_othery[0] ),
    .B(_03101_),
    .X(_03108_));
 sky130_fd_sc_hd__o211a_1 _19034_ (.A1(\rbzero.spi_registers.new_other[0] ),
    .A2(_03098_),
    .B1(_03108_),
    .C1(_03103_),
    .X(_00761_));
 sky130_fd_sc_hd__or2_1 _19035_ (.A(\rbzero.map_overlay.i_othery[1] ),
    .B(_03101_),
    .X(_03109_));
 sky130_fd_sc_hd__buf_6 _19036_ (.A(_08116_),
    .X(_03110_));
 sky130_fd_sc_hd__buf_2 _19037_ (.A(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__o211a_1 _19038_ (.A1(\rbzero.spi_registers.new_other[1] ),
    .A2(_03098_),
    .B1(_03109_),
    .C1(_03111_),
    .X(_00762_));
 sky130_fd_sc_hd__or2_1 _19039_ (.A(\rbzero.map_overlay.i_othery[2] ),
    .B(_03101_),
    .X(_03112_));
 sky130_fd_sc_hd__o211a_1 _19040_ (.A1(\rbzero.spi_registers.new_other[2] ),
    .A2(_03098_),
    .B1(_03112_),
    .C1(_03111_),
    .X(_00763_));
 sky130_fd_sc_hd__or2_1 _19041_ (.A(\rbzero.map_overlay.i_othery[3] ),
    .B(_03101_),
    .X(_03113_));
 sky130_fd_sc_hd__o211a_1 _19042_ (.A1(\rbzero.spi_registers.new_other[3] ),
    .A2(_03098_),
    .B1(_03113_),
    .C1(_03111_),
    .X(_00764_));
 sky130_fd_sc_hd__or2_1 _19043_ (.A(\rbzero.map_overlay.i_othery[4] ),
    .B(_03101_),
    .X(_03114_));
 sky130_fd_sc_hd__o211a_1 _19044_ (.A1(\rbzero.spi_registers.new_other[4] ),
    .A2(_03098_),
    .B1(_03114_),
    .C1(_03111_),
    .X(_00765_));
 sky130_fd_sc_hd__inv_2 _19045_ (.A(\rbzero.spi_registers.got_new_vinf ),
    .Y(_03115_));
 sky130_fd_sc_hd__nand3_4 _19046_ (.A(_05270_),
    .B(_03091_),
    .C(_03093_),
    .Y(_03116_));
 sky130_fd_sc_hd__a21o_1 _19047_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_03100_),
    .B1(\rbzero.row_render.vinf ),
    .X(_03117_));
 sky130_fd_sc_hd__clkbuf_8 _19048_ (.A(_03084_),
    .X(_03118_));
 sky130_fd_sc_hd__o311a_1 _19049_ (.A1(\rbzero.spi_registers.new_vinf ),
    .A2(_03115_),
    .A3(_03116_),
    .B1(_03117_),
    .C1(_03118_),
    .X(_00766_));
 sky130_fd_sc_hd__nand2_2 _19050_ (.A(\rbzero.spi_registers.got_new_mapd ),
    .B(_03096_),
    .Y(_03119_));
 sky130_fd_sc_hd__buf_2 _19051_ (.A(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__and2_1 _19052_ (.A(\rbzero.spi_registers.got_new_mapd ),
    .B(_03100_),
    .X(_03121_));
 sky130_fd_sc_hd__clkbuf_2 _19053_ (.A(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__or2_1 _19054_ (.A(\rbzero.map_overlay.i_mapdx[0] ),
    .B(_03122_),
    .X(_03123_));
 sky130_fd_sc_hd__o211a_1 _19055_ (.A1(\rbzero.spi_registers.new_mapd[10] ),
    .A2(_03120_),
    .B1(_03123_),
    .C1(_03111_),
    .X(_00767_));
 sky130_fd_sc_hd__or2_1 _19056_ (.A(\rbzero.map_overlay.i_mapdx[1] ),
    .B(_03122_),
    .X(_03124_));
 sky130_fd_sc_hd__o211a_1 _19057_ (.A1(\rbzero.spi_registers.new_mapd[11] ),
    .A2(_03120_),
    .B1(_03124_),
    .C1(_03111_),
    .X(_00768_));
 sky130_fd_sc_hd__or2_1 _19058_ (.A(\rbzero.map_overlay.i_mapdx[2] ),
    .B(_03122_),
    .X(_03125_));
 sky130_fd_sc_hd__o211a_1 _19059_ (.A1(\rbzero.spi_registers.new_mapd[12] ),
    .A2(_03120_),
    .B1(_03125_),
    .C1(_03111_),
    .X(_00769_));
 sky130_fd_sc_hd__or2_1 _19060_ (.A(\rbzero.map_overlay.i_mapdx[3] ),
    .B(_03122_),
    .X(_03126_));
 sky130_fd_sc_hd__o211a_1 _19061_ (.A1(\rbzero.spi_registers.new_mapd[13] ),
    .A2(_03120_),
    .B1(_03126_),
    .C1(_03111_),
    .X(_00770_));
 sky130_fd_sc_hd__or2_1 _19062_ (.A(\rbzero.map_overlay.i_mapdx[4] ),
    .B(_03122_),
    .X(_03127_));
 sky130_fd_sc_hd__o211a_1 _19063_ (.A1(\rbzero.spi_registers.new_mapd[14] ),
    .A2(_03120_),
    .B1(_03127_),
    .C1(_03111_),
    .X(_00771_));
 sky130_fd_sc_hd__or2_1 _19064_ (.A(\rbzero.map_overlay.i_mapdx[5] ),
    .B(_03122_),
    .X(_03128_));
 sky130_fd_sc_hd__o211a_1 _19065_ (.A1(\rbzero.spi_registers.new_mapd[15] ),
    .A2(_03120_),
    .B1(_03128_),
    .C1(_03111_),
    .X(_00772_));
 sky130_fd_sc_hd__or2_1 _19066_ (.A(\rbzero.map_overlay.i_mapdy[0] ),
    .B(_03122_),
    .X(_03129_));
 sky130_fd_sc_hd__buf_2 _19067_ (.A(_03110_),
    .X(_03130_));
 sky130_fd_sc_hd__o211a_1 _19068_ (.A1(\rbzero.spi_registers.new_mapd[4] ),
    .A2(_03120_),
    .B1(_03129_),
    .C1(_03130_),
    .X(_00773_));
 sky130_fd_sc_hd__or2_1 _19069_ (.A(\rbzero.map_overlay.i_mapdy[1] ),
    .B(_03122_),
    .X(_03131_));
 sky130_fd_sc_hd__o211a_1 _19070_ (.A1(\rbzero.spi_registers.new_mapd[5] ),
    .A2(_03120_),
    .B1(_03131_),
    .C1(_03130_),
    .X(_00774_));
 sky130_fd_sc_hd__or2_1 _19071_ (.A(\rbzero.map_overlay.i_mapdy[2] ),
    .B(_03122_),
    .X(_03132_));
 sky130_fd_sc_hd__o211a_1 _19072_ (.A1(\rbzero.spi_registers.new_mapd[6] ),
    .A2(_03120_),
    .B1(_03132_),
    .C1(_03130_),
    .X(_00775_));
 sky130_fd_sc_hd__or2_1 _19073_ (.A(\rbzero.map_overlay.i_mapdy[3] ),
    .B(_03122_),
    .X(_03133_));
 sky130_fd_sc_hd__o211a_1 _19074_ (.A1(\rbzero.spi_registers.new_mapd[7] ),
    .A2(_03120_),
    .B1(_03133_),
    .C1(_03130_),
    .X(_00776_));
 sky130_fd_sc_hd__or2_1 _19075_ (.A(\rbzero.map_overlay.i_mapdy[4] ),
    .B(_03121_),
    .X(_03134_));
 sky130_fd_sc_hd__o211a_1 _19076_ (.A1(\rbzero.spi_registers.new_mapd[8] ),
    .A2(_03119_),
    .B1(_03134_),
    .C1(_03130_),
    .X(_00777_));
 sky130_fd_sc_hd__or2_1 _19077_ (.A(\rbzero.map_overlay.i_mapdy[5] ),
    .B(_03121_),
    .X(_03135_));
 sky130_fd_sc_hd__o211a_1 _19078_ (.A1(\rbzero.spi_registers.new_mapd[9] ),
    .A2(_03119_),
    .B1(_03135_),
    .C1(_03130_),
    .X(_00778_));
 sky130_fd_sc_hd__or2_1 _19079_ (.A(\rbzero.mapdxw[0] ),
    .B(_03121_),
    .X(_03136_));
 sky130_fd_sc_hd__o211a_1 _19080_ (.A1(\rbzero.spi_registers.new_mapd[2] ),
    .A2(_03119_),
    .B1(_03136_),
    .C1(_03130_),
    .X(_00779_));
 sky130_fd_sc_hd__or2_1 _19081_ (.A(\rbzero.mapdxw[1] ),
    .B(_03121_),
    .X(_03137_));
 sky130_fd_sc_hd__o211a_1 _19082_ (.A1(\rbzero.spi_registers.new_mapd[3] ),
    .A2(_03119_),
    .B1(_03137_),
    .C1(_03130_),
    .X(_00780_));
 sky130_fd_sc_hd__or2_1 _19083_ (.A(\rbzero.mapdyw[0] ),
    .B(_03121_),
    .X(_03138_));
 sky130_fd_sc_hd__o211a_1 _19084_ (.A1(\rbzero.spi_registers.new_mapd[0] ),
    .A2(_03119_),
    .B1(_03138_),
    .C1(_03130_),
    .X(_00781_));
 sky130_fd_sc_hd__or2_1 _19085_ (.A(\rbzero.mapdyw[1] ),
    .B(_03121_),
    .X(_03139_));
 sky130_fd_sc_hd__o211a_1 _19086_ (.A1(\rbzero.spi_registers.new_mapd[1] ),
    .A2(_03119_),
    .B1(_03139_),
    .C1(_03130_),
    .X(_00782_));
 sky130_fd_sc_hd__nand2_2 _19087_ (.A(\rbzero.spi_registers.got_new_texadd[0] ),
    .B(_03096_),
    .Y(_03140_));
 sky130_fd_sc_hd__clkbuf_4 _19088_ (.A(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__and2_1 _19089_ (.A(\rbzero.spi_registers.got_new_texadd[0] ),
    .B(_03100_),
    .X(_03142_));
 sky130_fd_sc_hd__buf_2 _19090_ (.A(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__or2_1 _19091_ (.A(\rbzero.spi_registers.texadd0[0] ),
    .B(_03143_),
    .X(_03144_));
 sky130_fd_sc_hd__clkbuf_4 _19092_ (.A(_03110_),
    .X(_03145_));
 sky130_fd_sc_hd__o211a_1 _19093_ (.A1(\rbzero.spi_registers.new_texadd[0][0] ),
    .A2(_03141_),
    .B1(_03144_),
    .C1(_03145_),
    .X(_00783_));
 sky130_fd_sc_hd__or2_1 _19094_ (.A(\rbzero.spi_registers.texadd0[1] ),
    .B(_03143_),
    .X(_03146_));
 sky130_fd_sc_hd__o211a_1 _19095_ (.A1(\rbzero.spi_registers.new_texadd[0][1] ),
    .A2(_03141_),
    .B1(_03146_),
    .C1(_03145_),
    .X(_00784_));
 sky130_fd_sc_hd__or2_1 _19096_ (.A(\rbzero.spi_registers.texadd0[2] ),
    .B(_03143_),
    .X(_03147_));
 sky130_fd_sc_hd__o211a_1 _19097_ (.A1(\rbzero.spi_registers.new_texadd[0][2] ),
    .A2(_03141_),
    .B1(_03147_),
    .C1(_03145_),
    .X(_00785_));
 sky130_fd_sc_hd__or2_1 _19098_ (.A(\rbzero.spi_registers.texadd0[3] ),
    .B(_03143_),
    .X(_03148_));
 sky130_fd_sc_hd__o211a_1 _19099_ (.A1(\rbzero.spi_registers.new_texadd[0][3] ),
    .A2(_03141_),
    .B1(_03148_),
    .C1(_03145_),
    .X(_00786_));
 sky130_fd_sc_hd__or2_1 _19100_ (.A(\rbzero.spi_registers.texadd0[4] ),
    .B(_03143_),
    .X(_03149_));
 sky130_fd_sc_hd__o211a_1 _19101_ (.A1(\rbzero.spi_registers.new_texadd[0][4] ),
    .A2(_03141_),
    .B1(_03149_),
    .C1(_03145_),
    .X(_00787_));
 sky130_fd_sc_hd__or2_1 _19102_ (.A(\rbzero.spi_registers.texadd0[5] ),
    .B(_03143_),
    .X(_03150_));
 sky130_fd_sc_hd__o211a_1 _19103_ (.A1(\rbzero.spi_registers.new_texadd[0][5] ),
    .A2(_03141_),
    .B1(_03150_),
    .C1(_03145_),
    .X(_00788_));
 sky130_fd_sc_hd__or2_1 _19104_ (.A(\rbzero.spi_registers.texadd0[6] ),
    .B(_03143_),
    .X(_03151_));
 sky130_fd_sc_hd__o211a_1 _19105_ (.A1(\rbzero.spi_registers.new_texadd[0][6] ),
    .A2(_03141_),
    .B1(_03151_),
    .C1(_03145_),
    .X(_00789_));
 sky130_fd_sc_hd__or2_1 _19106_ (.A(\rbzero.spi_registers.texadd0[7] ),
    .B(_03143_),
    .X(_03152_));
 sky130_fd_sc_hd__o211a_1 _19107_ (.A1(\rbzero.spi_registers.new_texadd[0][7] ),
    .A2(_03141_),
    .B1(_03152_),
    .C1(_03145_),
    .X(_00790_));
 sky130_fd_sc_hd__or2_1 _19108_ (.A(\rbzero.spi_registers.texadd0[8] ),
    .B(_03143_),
    .X(_03153_));
 sky130_fd_sc_hd__o211a_1 _19109_ (.A1(\rbzero.spi_registers.new_texadd[0][8] ),
    .A2(_03141_),
    .B1(_03153_),
    .C1(_03145_),
    .X(_00791_));
 sky130_fd_sc_hd__or2_1 _19110_ (.A(\rbzero.spi_registers.texadd0[9] ),
    .B(_03143_),
    .X(_03154_));
 sky130_fd_sc_hd__o211a_1 _19111_ (.A1(\rbzero.spi_registers.new_texadd[0][9] ),
    .A2(_03141_),
    .B1(_03154_),
    .C1(_03145_),
    .X(_00792_));
 sky130_fd_sc_hd__clkbuf_4 _19112_ (.A(_03140_),
    .X(_03155_));
 sky130_fd_sc_hd__clkbuf_2 _19113_ (.A(_03142_),
    .X(_03156_));
 sky130_fd_sc_hd__or2_1 _19114_ (.A(\rbzero.spi_registers.texadd0[10] ),
    .B(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__clkbuf_4 _19115_ (.A(_03110_),
    .X(_03158_));
 sky130_fd_sc_hd__o211a_1 _19116_ (.A1(\rbzero.spi_registers.new_texadd[0][10] ),
    .A2(_03155_),
    .B1(_03157_),
    .C1(_03158_),
    .X(_00793_));
 sky130_fd_sc_hd__or2_1 _19117_ (.A(\rbzero.spi_registers.texadd0[11] ),
    .B(_03156_),
    .X(_03159_));
 sky130_fd_sc_hd__o211a_1 _19118_ (.A1(\rbzero.spi_registers.new_texadd[0][11] ),
    .A2(_03155_),
    .B1(_03159_),
    .C1(_03158_),
    .X(_00794_));
 sky130_fd_sc_hd__or2_1 _19119_ (.A(\rbzero.spi_registers.texadd0[12] ),
    .B(_03156_),
    .X(_03160_));
 sky130_fd_sc_hd__o211a_1 _19120_ (.A1(\rbzero.spi_registers.new_texadd[0][12] ),
    .A2(_03155_),
    .B1(_03160_),
    .C1(_03158_),
    .X(_00795_));
 sky130_fd_sc_hd__or2_1 _19121_ (.A(\rbzero.spi_registers.texadd0[13] ),
    .B(_03156_),
    .X(_03161_));
 sky130_fd_sc_hd__o211a_1 _19122_ (.A1(\rbzero.spi_registers.new_texadd[0][13] ),
    .A2(_03155_),
    .B1(_03161_),
    .C1(_03158_),
    .X(_00796_));
 sky130_fd_sc_hd__or2_1 _19123_ (.A(\rbzero.spi_registers.texadd0[14] ),
    .B(_03156_),
    .X(_03162_));
 sky130_fd_sc_hd__o211a_1 _19124_ (.A1(\rbzero.spi_registers.new_texadd[0][14] ),
    .A2(_03155_),
    .B1(_03162_),
    .C1(_03158_),
    .X(_00797_));
 sky130_fd_sc_hd__or2_1 _19125_ (.A(\rbzero.spi_registers.texadd0[15] ),
    .B(_03156_),
    .X(_03163_));
 sky130_fd_sc_hd__o211a_1 _19126_ (.A1(\rbzero.spi_registers.new_texadd[0][15] ),
    .A2(_03155_),
    .B1(_03163_),
    .C1(_03158_),
    .X(_00798_));
 sky130_fd_sc_hd__or2_1 _19127_ (.A(\rbzero.spi_registers.texadd0[16] ),
    .B(_03156_),
    .X(_03164_));
 sky130_fd_sc_hd__o211a_1 _19128_ (.A1(\rbzero.spi_registers.new_texadd[0][16] ),
    .A2(_03155_),
    .B1(_03164_),
    .C1(_03158_),
    .X(_00799_));
 sky130_fd_sc_hd__or2_1 _19129_ (.A(\rbzero.spi_registers.texadd0[17] ),
    .B(_03156_),
    .X(_03165_));
 sky130_fd_sc_hd__o211a_1 _19130_ (.A1(\rbzero.spi_registers.new_texadd[0][17] ),
    .A2(_03155_),
    .B1(_03165_),
    .C1(_03158_),
    .X(_00800_));
 sky130_fd_sc_hd__or2_1 _19131_ (.A(\rbzero.spi_registers.texadd0[18] ),
    .B(_03156_),
    .X(_03166_));
 sky130_fd_sc_hd__o211a_1 _19132_ (.A1(\rbzero.spi_registers.new_texadd[0][18] ),
    .A2(_03155_),
    .B1(_03166_),
    .C1(_03158_),
    .X(_00801_));
 sky130_fd_sc_hd__or2_1 _19133_ (.A(\rbzero.spi_registers.texadd0[19] ),
    .B(_03156_),
    .X(_03167_));
 sky130_fd_sc_hd__o211a_1 _19134_ (.A1(\rbzero.spi_registers.new_texadd[0][19] ),
    .A2(_03155_),
    .B1(_03167_),
    .C1(_03158_),
    .X(_00802_));
 sky130_fd_sc_hd__or2_1 _19135_ (.A(\rbzero.spi_registers.texadd0[20] ),
    .B(_03142_),
    .X(_03168_));
 sky130_fd_sc_hd__clkbuf_4 _19136_ (.A(_03110_),
    .X(_03169_));
 sky130_fd_sc_hd__o211a_1 _19137_ (.A1(\rbzero.spi_registers.new_texadd[0][20] ),
    .A2(_03140_),
    .B1(_03168_),
    .C1(_03169_),
    .X(_00803_));
 sky130_fd_sc_hd__or2_1 _19138_ (.A(\rbzero.spi_registers.texadd0[21] ),
    .B(_03142_),
    .X(_03170_));
 sky130_fd_sc_hd__o211a_1 _19139_ (.A1(\rbzero.spi_registers.new_texadd[0][21] ),
    .A2(_03140_),
    .B1(_03170_),
    .C1(_03169_),
    .X(_00804_));
 sky130_fd_sc_hd__or2_1 _19140_ (.A(\rbzero.spi_registers.texadd0[22] ),
    .B(_03142_),
    .X(_03171_));
 sky130_fd_sc_hd__o211a_1 _19141_ (.A1(\rbzero.spi_registers.new_texadd[0][22] ),
    .A2(_03140_),
    .B1(_03171_),
    .C1(_03169_),
    .X(_00805_));
 sky130_fd_sc_hd__or2_1 _19142_ (.A(\rbzero.spi_registers.texadd0[23] ),
    .B(_03142_),
    .X(_03172_));
 sky130_fd_sc_hd__o211a_1 _19143_ (.A1(\rbzero.spi_registers.new_texadd[0][23] ),
    .A2(_03140_),
    .B1(_03172_),
    .C1(_03169_),
    .X(_00806_));
 sky130_fd_sc_hd__nand2_2 _19144_ (.A(\rbzero.spi_registers.got_new_texadd[1] ),
    .B(_03096_),
    .Y(_03173_));
 sky130_fd_sc_hd__clkbuf_4 _19145_ (.A(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__and2_1 _19146_ (.A(\rbzero.spi_registers.got_new_texadd[1] ),
    .B(_03100_),
    .X(_03175_));
 sky130_fd_sc_hd__buf_2 _19147_ (.A(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__or2_1 _19148_ (.A(\rbzero.spi_registers.texadd1[0] ),
    .B(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__o211a_1 _19149_ (.A1(\rbzero.spi_registers.new_texadd[1][0] ),
    .A2(_03174_),
    .B1(_03177_),
    .C1(_03169_),
    .X(_00807_));
 sky130_fd_sc_hd__or2_1 _19150_ (.A(\rbzero.spi_registers.texadd1[1] ),
    .B(_03176_),
    .X(_03178_));
 sky130_fd_sc_hd__o211a_1 _19151_ (.A1(\rbzero.spi_registers.new_texadd[1][1] ),
    .A2(_03174_),
    .B1(_03178_),
    .C1(_03169_),
    .X(_00808_));
 sky130_fd_sc_hd__or2_1 _19152_ (.A(\rbzero.spi_registers.texadd1[2] ),
    .B(_03176_),
    .X(_03179_));
 sky130_fd_sc_hd__o211a_1 _19153_ (.A1(\rbzero.spi_registers.new_texadd[1][2] ),
    .A2(_03174_),
    .B1(_03179_),
    .C1(_03169_),
    .X(_00809_));
 sky130_fd_sc_hd__or2_1 _19154_ (.A(\rbzero.spi_registers.texadd1[3] ),
    .B(_03176_),
    .X(_03180_));
 sky130_fd_sc_hd__o211a_1 _19155_ (.A1(\rbzero.spi_registers.new_texadd[1][3] ),
    .A2(_03174_),
    .B1(_03180_),
    .C1(_03169_),
    .X(_00810_));
 sky130_fd_sc_hd__or2_1 _19156_ (.A(\rbzero.spi_registers.texadd1[4] ),
    .B(_03176_),
    .X(_03181_));
 sky130_fd_sc_hd__o211a_1 _19157_ (.A1(\rbzero.spi_registers.new_texadd[1][4] ),
    .A2(_03174_),
    .B1(_03181_),
    .C1(_03169_),
    .X(_00811_));
 sky130_fd_sc_hd__or2_1 _19158_ (.A(\rbzero.spi_registers.texadd1[5] ),
    .B(_03176_),
    .X(_03182_));
 sky130_fd_sc_hd__o211a_1 _19159_ (.A1(\rbzero.spi_registers.new_texadd[1][5] ),
    .A2(_03174_),
    .B1(_03182_),
    .C1(_03169_),
    .X(_00812_));
 sky130_fd_sc_hd__or2_1 _19160_ (.A(\rbzero.spi_registers.texadd1[6] ),
    .B(_03176_),
    .X(_03183_));
 sky130_fd_sc_hd__clkbuf_4 _19161_ (.A(_03110_),
    .X(_03184_));
 sky130_fd_sc_hd__o211a_1 _19162_ (.A1(\rbzero.spi_registers.new_texadd[1][6] ),
    .A2(_03174_),
    .B1(_03183_),
    .C1(_03184_),
    .X(_00813_));
 sky130_fd_sc_hd__or2_1 _19163_ (.A(\rbzero.spi_registers.texadd1[7] ),
    .B(_03176_),
    .X(_03185_));
 sky130_fd_sc_hd__o211a_1 _19164_ (.A1(\rbzero.spi_registers.new_texadd[1][7] ),
    .A2(_03174_),
    .B1(_03185_),
    .C1(_03184_),
    .X(_00814_));
 sky130_fd_sc_hd__or2_1 _19165_ (.A(\rbzero.spi_registers.texadd1[8] ),
    .B(_03176_),
    .X(_03186_));
 sky130_fd_sc_hd__o211a_1 _19166_ (.A1(\rbzero.spi_registers.new_texadd[1][8] ),
    .A2(_03174_),
    .B1(_03186_),
    .C1(_03184_),
    .X(_00815_));
 sky130_fd_sc_hd__or2_1 _19167_ (.A(\rbzero.spi_registers.texadd1[9] ),
    .B(_03176_),
    .X(_03187_));
 sky130_fd_sc_hd__o211a_1 _19168_ (.A1(\rbzero.spi_registers.new_texadd[1][9] ),
    .A2(_03174_),
    .B1(_03187_),
    .C1(_03184_),
    .X(_00816_));
 sky130_fd_sc_hd__clkbuf_4 _19169_ (.A(_03173_),
    .X(_03188_));
 sky130_fd_sc_hd__buf_2 _19170_ (.A(_03175_),
    .X(_03189_));
 sky130_fd_sc_hd__or2_1 _19171_ (.A(\rbzero.spi_registers.texadd1[10] ),
    .B(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__o211a_1 _19172_ (.A1(\rbzero.spi_registers.new_texadd[1][10] ),
    .A2(_03188_),
    .B1(_03190_),
    .C1(_03184_),
    .X(_00817_));
 sky130_fd_sc_hd__or2_1 _19173_ (.A(\rbzero.spi_registers.texadd1[11] ),
    .B(_03189_),
    .X(_03191_));
 sky130_fd_sc_hd__o211a_1 _19174_ (.A1(\rbzero.spi_registers.new_texadd[1][11] ),
    .A2(_03188_),
    .B1(_03191_),
    .C1(_03184_),
    .X(_00818_));
 sky130_fd_sc_hd__or2_1 _19175_ (.A(\rbzero.spi_registers.texadd1[12] ),
    .B(_03189_),
    .X(_03192_));
 sky130_fd_sc_hd__o211a_1 _19176_ (.A1(\rbzero.spi_registers.new_texadd[1][12] ),
    .A2(_03188_),
    .B1(_03192_),
    .C1(_03184_),
    .X(_00819_));
 sky130_fd_sc_hd__or2_1 _19177_ (.A(\rbzero.spi_registers.texadd1[13] ),
    .B(_03189_),
    .X(_03193_));
 sky130_fd_sc_hd__o211a_1 _19178_ (.A1(\rbzero.spi_registers.new_texadd[1][13] ),
    .A2(_03188_),
    .B1(_03193_),
    .C1(_03184_),
    .X(_00820_));
 sky130_fd_sc_hd__or2_1 _19179_ (.A(\rbzero.spi_registers.texadd1[14] ),
    .B(_03189_),
    .X(_03194_));
 sky130_fd_sc_hd__o211a_1 _19180_ (.A1(\rbzero.spi_registers.new_texadd[1][14] ),
    .A2(_03188_),
    .B1(_03194_),
    .C1(_03184_),
    .X(_00821_));
 sky130_fd_sc_hd__or2_1 _19181_ (.A(\rbzero.spi_registers.texadd1[15] ),
    .B(_03189_),
    .X(_03195_));
 sky130_fd_sc_hd__o211a_1 _19182_ (.A1(\rbzero.spi_registers.new_texadd[1][15] ),
    .A2(_03188_),
    .B1(_03195_),
    .C1(_03184_),
    .X(_00822_));
 sky130_fd_sc_hd__or2_1 _19183_ (.A(\rbzero.spi_registers.texadd1[16] ),
    .B(_03189_),
    .X(_03196_));
 sky130_fd_sc_hd__clkbuf_4 _19184_ (.A(_03110_),
    .X(_03197_));
 sky130_fd_sc_hd__o211a_1 _19185_ (.A1(\rbzero.spi_registers.new_texadd[1][16] ),
    .A2(_03188_),
    .B1(_03196_),
    .C1(_03197_),
    .X(_00823_));
 sky130_fd_sc_hd__or2_1 _19186_ (.A(\rbzero.spi_registers.texadd1[17] ),
    .B(_03189_),
    .X(_03198_));
 sky130_fd_sc_hd__o211a_1 _19187_ (.A1(\rbzero.spi_registers.new_texadd[1][17] ),
    .A2(_03188_),
    .B1(_03198_),
    .C1(_03197_),
    .X(_00824_));
 sky130_fd_sc_hd__or2_1 _19188_ (.A(\rbzero.spi_registers.texadd1[18] ),
    .B(_03189_),
    .X(_03199_));
 sky130_fd_sc_hd__o211a_1 _19189_ (.A1(\rbzero.spi_registers.new_texadd[1][18] ),
    .A2(_03188_),
    .B1(_03199_),
    .C1(_03197_),
    .X(_00825_));
 sky130_fd_sc_hd__or2_1 _19190_ (.A(\rbzero.spi_registers.texadd1[19] ),
    .B(_03189_),
    .X(_03200_));
 sky130_fd_sc_hd__o211a_1 _19191_ (.A1(\rbzero.spi_registers.new_texadd[1][19] ),
    .A2(_03188_),
    .B1(_03200_),
    .C1(_03197_),
    .X(_00826_));
 sky130_fd_sc_hd__or2_1 _19192_ (.A(\rbzero.spi_registers.texadd1[20] ),
    .B(_03175_),
    .X(_03201_));
 sky130_fd_sc_hd__o211a_1 _19193_ (.A1(\rbzero.spi_registers.new_texadd[1][20] ),
    .A2(_03173_),
    .B1(_03201_),
    .C1(_03197_),
    .X(_00827_));
 sky130_fd_sc_hd__or2_1 _19194_ (.A(\rbzero.spi_registers.texadd1[21] ),
    .B(_03175_),
    .X(_03202_));
 sky130_fd_sc_hd__o211a_1 _19195_ (.A1(\rbzero.spi_registers.new_texadd[1][21] ),
    .A2(_03173_),
    .B1(_03202_),
    .C1(_03197_),
    .X(_00828_));
 sky130_fd_sc_hd__or2_1 _19196_ (.A(\rbzero.spi_registers.texadd1[22] ),
    .B(_03175_),
    .X(_03203_));
 sky130_fd_sc_hd__o211a_1 _19197_ (.A1(\rbzero.spi_registers.new_texadd[1][22] ),
    .A2(_03173_),
    .B1(_03203_),
    .C1(_03197_),
    .X(_00829_));
 sky130_fd_sc_hd__or2_1 _19198_ (.A(\rbzero.spi_registers.texadd1[23] ),
    .B(_03175_),
    .X(_03204_));
 sky130_fd_sc_hd__o211a_1 _19199_ (.A1(\rbzero.spi_registers.new_texadd[1][23] ),
    .A2(_03173_),
    .B1(_03204_),
    .C1(_03197_),
    .X(_00830_));
 sky130_fd_sc_hd__nand2_2 _19200_ (.A(\rbzero.spi_registers.got_new_texadd[2] ),
    .B(_03096_),
    .Y(_03205_));
 sky130_fd_sc_hd__clkbuf_4 _19201_ (.A(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__and2_2 _19202_ (.A(\rbzero.spi_registers.got_new_texadd[2] ),
    .B(_03100_),
    .X(_03207_));
 sky130_fd_sc_hd__buf_2 _19203_ (.A(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__or2_1 _19204_ (.A(\rbzero.spi_registers.texadd2[0] ),
    .B(_03208_),
    .X(_03209_));
 sky130_fd_sc_hd__o211a_1 _19205_ (.A1(\rbzero.spi_registers.new_texadd[2][0] ),
    .A2(_03206_),
    .B1(_03209_),
    .C1(_03197_),
    .X(_00831_));
 sky130_fd_sc_hd__or2_1 _19206_ (.A(\rbzero.spi_registers.texadd2[1] ),
    .B(_03208_),
    .X(_03210_));
 sky130_fd_sc_hd__o211a_1 _19207_ (.A1(\rbzero.spi_registers.new_texadd[2][1] ),
    .A2(_03206_),
    .B1(_03210_),
    .C1(_03197_),
    .X(_00832_));
 sky130_fd_sc_hd__or2_1 _19208_ (.A(\rbzero.spi_registers.texadd2[2] ),
    .B(_03208_),
    .X(_03211_));
 sky130_fd_sc_hd__buf_6 _19209_ (.A(_08116_),
    .X(_03212_));
 sky130_fd_sc_hd__clkbuf_4 _19210_ (.A(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__o211a_1 _19211_ (.A1(\rbzero.spi_registers.new_texadd[2][2] ),
    .A2(_03206_),
    .B1(_03211_),
    .C1(_03213_),
    .X(_00833_));
 sky130_fd_sc_hd__or2_1 _19212_ (.A(\rbzero.spi_registers.texadd2[3] ),
    .B(_03208_),
    .X(_03214_));
 sky130_fd_sc_hd__o211a_1 _19213_ (.A1(\rbzero.spi_registers.new_texadd[2][3] ),
    .A2(_03206_),
    .B1(_03214_),
    .C1(_03213_),
    .X(_00834_));
 sky130_fd_sc_hd__or2_1 _19214_ (.A(\rbzero.spi_registers.texadd2[4] ),
    .B(_03208_),
    .X(_03215_));
 sky130_fd_sc_hd__o211a_1 _19215_ (.A1(\rbzero.spi_registers.new_texadd[2][4] ),
    .A2(_03206_),
    .B1(_03215_),
    .C1(_03213_),
    .X(_00835_));
 sky130_fd_sc_hd__or2_1 _19216_ (.A(\rbzero.spi_registers.texadd2[5] ),
    .B(_03208_),
    .X(_03216_));
 sky130_fd_sc_hd__o211a_1 _19217_ (.A1(\rbzero.spi_registers.new_texadd[2][5] ),
    .A2(_03206_),
    .B1(_03216_),
    .C1(_03213_),
    .X(_00836_));
 sky130_fd_sc_hd__or2_1 _19218_ (.A(\rbzero.spi_registers.texadd2[6] ),
    .B(_03208_),
    .X(_03217_));
 sky130_fd_sc_hd__o211a_1 _19219_ (.A1(\rbzero.spi_registers.new_texadd[2][6] ),
    .A2(_03206_),
    .B1(_03217_),
    .C1(_03213_),
    .X(_00837_));
 sky130_fd_sc_hd__or2_1 _19220_ (.A(\rbzero.spi_registers.texadd2[7] ),
    .B(_03208_),
    .X(_03218_));
 sky130_fd_sc_hd__o211a_1 _19221_ (.A1(\rbzero.spi_registers.new_texadd[2][7] ),
    .A2(_03206_),
    .B1(_03218_),
    .C1(_03213_),
    .X(_00838_));
 sky130_fd_sc_hd__or2_1 _19222_ (.A(\rbzero.spi_registers.texadd2[8] ),
    .B(_03208_),
    .X(_03219_));
 sky130_fd_sc_hd__o211a_1 _19223_ (.A1(\rbzero.spi_registers.new_texadd[2][8] ),
    .A2(_03206_),
    .B1(_03219_),
    .C1(_03213_),
    .X(_00839_));
 sky130_fd_sc_hd__or2_1 _19224_ (.A(\rbzero.spi_registers.texadd2[9] ),
    .B(_03208_),
    .X(_03220_));
 sky130_fd_sc_hd__o211a_1 _19225_ (.A1(\rbzero.spi_registers.new_texadd[2][9] ),
    .A2(_03206_),
    .B1(_03220_),
    .C1(_03213_),
    .X(_00840_));
 sky130_fd_sc_hd__clkbuf_4 _19226_ (.A(_03205_),
    .X(_03221_));
 sky130_fd_sc_hd__buf_2 _19227_ (.A(_03207_),
    .X(_03222_));
 sky130_fd_sc_hd__or2_1 _19228_ (.A(\rbzero.spi_registers.texadd2[10] ),
    .B(_03222_),
    .X(_03223_));
 sky130_fd_sc_hd__o211a_1 _19229_ (.A1(\rbzero.spi_registers.new_texadd[2][10] ),
    .A2(_03221_),
    .B1(_03223_),
    .C1(_03213_),
    .X(_00841_));
 sky130_fd_sc_hd__or2_1 _19230_ (.A(\rbzero.spi_registers.texadd2[11] ),
    .B(_03222_),
    .X(_03224_));
 sky130_fd_sc_hd__o211a_1 _19231_ (.A1(\rbzero.spi_registers.new_texadd[2][11] ),
    .A2(_03221_),
    .B1(_03224_),
    .C1(_03213_),
    .X(_00842_));
 sky130_fd_sc_hd__or2_1 _19232_ (.A(\rbzero.spi_registers.texadd2[12] ),
    .B(_03222_),
    .X(_03225_));
 sky130_fd_sc_hd__clkbuf_4 _19233_ (.A(_03212_),
    .X(_03226_));
 sky130_fd_sc_hd__o211a_1 _19234_ (.A1(\rbzero.spi_registers.new_texadd[2][12] ),
    .A2(_03221_),
    .B1(_03225_),
    .C1(_03226_),
    .X(_00843_));
 sky130_fd_sc_hd__or2_1 _19235_ (.A(\rbzero.spi_registers.texadd2[13] ),
    .B(_03222_),
    .X(_03227_));
 sky130_fd_sc_hd__o211a_1 _19236_ (.A1(\rbzero.spi_registers.new_texadd[2][13] ),
    .A2(_03221_),
    .B1(_03227_),
    .C1(_03226_),
    .X(_00844_));
 sky130_fd_sc_hd__or2_1 _19237_ (.A(\rbzero.spi_registers.texadd2[14] ),
    .B(_03222_),
    .X(_03228_));
 sky130_fd_sc_hd__o211a_1 _19238_ (.A1(\rbzero.spi_registers.new_texadd[2][14] ),
    .A2(_03221_),
    .B1(_03228_),
    .C1(_03226_),
    .X(_00845_));
 sky130_fd_sc_hd__or2_1 _19239_ (.A(\rbzero.spi_registers.texadd2[15] ),
    .B(_03222_),
    .X(_03229_));
 sky130_fd_sc_hd__o211a_1 _19240_ (.A1(\rbzero.spi_registers.new_texadd[2][15] ),
    .A2(_03221_),
    .B1(_03229_),
    .C1(_03226_),
    .X(_00846_));
 sky130_fd_sc_hd__or2_1 _19241_ (.A(\rbzero.spi_registers.texadd2[16] ),
    .B(_03222_),
    .X(_03230_));
 sky130_fd_sc_hd__o211a_1 _19242_ (.A1(\rbzero.spi_registers.new_texadd[2][16] ),
    .A2(_03221_),
    .B1(_03230_),
    .C1(_03226_),
    .X(_00847_));
 sky130_fd_sc_hd__or2_1 _19243_ (.A(\rbzero.spi_registers.texadd2[17] ),
    .B(_03222_),
    .X(_03231_));
 sky130_fd_sc_hd__o211a_1 _19244_ (.A1(\rbzero.spi_registers.new_texadd[2][17] ),
    .A2(_03221_),
    .B1(_03231_),
    .C1(_03226_),
    .X(_00848_));
 sky130_fd_sc_hd__or2_1 _19245_ (.A(\rbzero.spi_registers.texadd2[18] ),
    .B(_03222_),
    .X(_03232_));
 sky130_fd_sc_hd__o211a_1 _19246_ (.A1(\rbzero.spi_registers.new_texadd[2][18] ),
    .A2(_03221_),
    .B1(_03232_),
    .C1(_03226_),
    .X(_00849_));
 sky130_fd_sc_hd__or2_1 _19247_ (.A(\rbzero.spi_registers.texadd2[19] ),
    .B(_03222_),
    .X(_03233_));
 sky130_fd_sc_hd__o211a_1 _19248_ (.A1(\rbzero.spi_registers.new_texadd[2][19] ),
    .A2(_03221_),
    .B1(_03233_),
    .C1(_03226_),
    .X(_00850_));
 sky130_fd_sc_hd__or2_1 _19249_ (.A(\rbzero.spi_registers.texadd2[20] ),
    .B(_03207_),
    .X(_03234_));
 sky130_fd_sc_hd__o211a_1 _19250_ (.A1(\rbzero.spi_registers.new_texadd[2][20] ),
    .A2(_03205_),
    .B1(_03234_),
    .C1(_03226_),
    .X(_00851_));
 sky130_fd_sc_hd__or2_1 _19251_ (.A(\rbzero.spi_registers.texadd2[21] ),
    .B(_03207_),
    .X(_03235_));
 sky130_fd_sc_hd__o211a_1 _19252_ (.A1(\rbzero.spi_registers.new_texadd[2][21] ),
    .A2(_03205_),
    .B1(_03235_),
    .C1(_03226_),
    .X(_00852_));
 sky130_fd_sc_hd__or2_1 _19253_ (.A(\rbzero.spi_registers.texadd2[22] ),
    .B(_03207_),
    .X(_03236_));
 sky130_fd_sc_hd__clkbuf_4 _19254_ (.A(_03212_),
    .X(_03237_));
 sky130_fd_sc_hd__o211a_1 _19255_ (.A1(\rbzero.spi_registers.new_texadd[2][22] ),
    .A2(_03205_),
    .B1(_03236_),
    .C1(_03237_),
    .X(_00853_));
 sky130_fd_sc_hd__or2_1 _19256_ (.A(\rbzero.spi_registers.texadd2[23] ),
    .B(_03207_),
    .X(_03238_));
 sky130_fd_sc_hd__o211a_1 _19257_ (.A1(\rbzero.spi_registers.new_texadd[2][23] ),
    .A2(_03205_),
    .B1(_03238_),
    .C1(_03237_),
    .X(_00854_));
 sky130_fd_sc_hd__nand2_2 _19258_ (.A(\rbzero.spi_registers.got_new_texadd[3] ),
    .B(_03096_),
    .Y(_03239_));
 sky130_fd_sc_hd__clkbuf_4 _19259_ (.A(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__and2_1 _19260_ (.A(\rbzero.spi_registers.got_new_texadd[3] ),
    .B(_03100_),
    .X(_03241_));
 sky130_fd_sc_hd__clkbuf_4 _19261_ (.A(_03241_),
    .X(_03242_));
 sky130_fd_sc_hd__or2_1 _19262_ (.A(\rbzero.spi_registers.texadd3[0] ),
    .B(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__o211a_1 _19263_ (.A1(\rbzero.spi_registers.new_texadd[3][0] ),
    .A2(_03240_),
    .B1(_03243_),
    .C1(_03237_),
    .X(_00855_));
 sky130_fd_sc_hd__or2_1 _19264_ (.A(\rbzero.spi_registers.texadd3[1] ),
    .B(_03242_),
    .X(_03244_));
 sky130_fd_sc_hd__o211a_1 _19265_ (.A1(\rbzero.spi_registers.new_texadd[3][1] ),
    .A2(_03240_),
    .B1(_03244_),
    .C1(_03237_),
    .X(_00856_));
 sky130_fd_sc_hd__or2_1 _19266_ (.A(\rbzero.spi_registers.texadd3[2] ),
    .B(_03242_),
    .X(_03245_));
 sky130_fd_sc_hd__o211a_1 _19267_ (.A1(\rbzero.spi_registers.new_texadd[3][2] ),
    .A2(_03240_),
    .B1(_03245_),
    .C1(_03237_),
    .X(_00857_));
 sky130_fd_sc_hd__or2_1 _19268_ (.A(\rbzero.spi_registers.texadd3[3] ),
    .B(_03242_),
    .X(_03246_));
 sky130_fd_sc_hd__o211a_1 _19269_ (.A1(\rbzero.spi_registers.new_texadd[3][3] ),
    .A2(_03240_),
    .B1(_03246_),
    .C1(_03237_),
    .X(_00858_));
 sky130_fd_sc_hd__or2_1 _19270_ (.A(\rbzero.spi_registers.texadd3[4] ),
    .B(_03242_),
    .X(_03247_));
 sky130_fd_sc_hd__o211a_1 _19271_ (.A1(\rbzero.spi_registers.new_texadd[3][4] ),
    .A2(_03240_),
    .B1(_03247_),
    .C1(_03237_),
    .X(_00859_));
 sky130_fd_sc_hd__or2_1 _19272_ (.A(\rbzero.spi_registers.texadd3[5] ),
    .B(_03242_),
    .X(_03248_));
 sky130_fd_sc_hd__o211a_1 _19273_ (.A1(\rbzero.spi_registers.new_texadd[3][5] ),
    .A2(_03240_),
    .B1(_03248_),
    .C1(_03237_),
    .X(_00860_));
 sky130_fd_sc_hd__or2_1 _19274_ (.A(\rbzero.spi_registers.texadd3[6] ),
    .B(_03242_),
    .X(_03249_));
 sky130_fd_sc_hd__o211a_1 _19275_ (.A1(\rbzero.spi_registers.new_texadd[3][6] ),
    .A2(_03240_),
    .B1(_03249_),
    .C1(_03237_),
    .X(_00861_));
 sky130_fd_sc_hd__or2_1 _19276_ (.A(\rbzero.spi_registers.texadd3[7] ),
    .B(_03242_),
    .X(_03250_));
 sky130_fd_sc_hd__o211a_1 _19277_ (.A1(\rbzero.spi_registers.new_texadd[3][7] ),
    .A2(_03240_),
    .B1(_03250_),
    .C1(_03237_),
    .X(_00862_));
 sky130_fd_sc_hd__or2_1 _19278_ (.A(\rbzero.spi_registers.texadd3[8] ),
    .B(_03242_),
    .X(_03251_));
 sky130_fd_sc_hd__clkbuf_4 _19279_ (.A(_03212_),
    .X(_03252_));
 sky130_fd_sc_hd__o211a_1 _19280_ (.A1(\rbzero.spi_registers.new_texadd[3][8] ),
    .A2(_03240_),
    .B1(_03251_),
    .C1(_03252_),
    .X(_00863_));
 sky130_fd_sc_hd__or2_1 _19281_ (.A(\rbzero.spi_registers.texadd3[9] ),
    .B(_03242_),
    .X(_03253_));
 sky130_fd_sc_hd__o211a_1 _19282_ (.A1(\rbzero.spi_registers.new_texadd[3][9] ),
    .A2(_03240_),
    .B1(_03253_),
    .C1(_03252_),
    .X(_00864_));
 sky130_fd_sc_hd__clkbuf_4 _19283_ (.A(_03239_),
    .X(_03254_));
 sky130_fd_sc_hd__buf_2 _19284_ (.A(_03241_),
    .X(_03255_));
 sky130_fd_sc_hd__or2_1 _19285_ (.A(\rbzero.spi_registers.texadd3[10] ),
    .B(_03255_),
    .X(_03256_));
 sky130_fd_sc_hd__o211a_1 _19286_ (.A1(\rbzero.spi_registers.new_texadd[3][10] ),
    .A2(_03254_),
    .B1(_03256_),
    .C1(_03252_),
    .X(_00865_));
 sky130_fd_sc_hd__or2_1 _19287_ (.A(\rbzero.spi_registers.texadd3[11] ),
    .B(_03255_),
    .X(_03257_));
 sky130_fd_sc_hd__o211a_1 _19288_ (.A1(\rbzero.spi_registers.new_texadd[3][11] ),
    .A2(_03254_),
    .B1(_03257_),
    .C1(_03252_),
    .X(_00866_));
 sky130_fd_sc_hd__or2_1 _19289_ (.A(\rbzero.spi_registers.texadd3[12] ),
    .B(_03255_),
    .X(_03258_));
 sky130_fd_sc_hd__o211a_1 _19290_ (.A1(\rbzero.spi_registers.new_texadd[3][12] ),
    .A2(_03254_),
    .B1(_03258_),
    .C1(_03252_),
    .X(_00867_));
 sky130_fd_sc_hd__or2_1 _19291_ (.A(\rbzero.spi_registers.texadd3[13] ),
    .B(_03255_),
    .X(_03259_));
 sky130_fd_sc_hd__o211a_1 _19292_ (.A1(\rbzero.spi_registers.new_texadd[3][13] ),
    .A2(_03254_),
    .B1(_03259_),
    .C1(_03252_),
    .X(_00868_));
 sky130_fd_sc_hd__or2_1 _19293_ (.A(\rbzero.spi_registers.texadd3[14] ),
    .B(_03255_),
    .X(_03260_));
 sky130_fd_sc_hd__o211a_1 _19294_ (.A1(\rbzero.spi_registers.new_texadd[3][14] ),
    .A2(_03254_),
    .B1(_03260_),
    .C1(_03252_),
    .X(_00869_));
 sky130_fd_sc_hd__or2_1 _19295_ (.A(\rbzero.spi_registers.texadd3[15] ),
    .B(_03255_),
    .X(_03261_));
 sky130_fd_sc_hd__o211a_1 _19296_ (.A1(\rbzero.spi_registers.new_texadd[3][15] ),
    .A2(_03254_),
    .B1(_03261_),
    .C1(_03252_),
    .X(_00870_));
 sky130_fd_sc_hd__or2_1 _19297_ (.A(\rbzero.spi_registers.texadd3[16] ),
    .B(_03255_),
    .X(_03262_));
 sky130_fd_sc_hd__o211a_1 _19298_ (.A1(\rbzero.spi_registers.new_texadd[3][16] ),
    .A2(_03254_),
    .B1(_03262_),
    .C1(_03252_),
    .X(_00871_));
 sky130_fd_sc_hd__or2_1 _19299_ (.A(\rbzero.spi_registers.texadd3[17] ),
    .B(_03255_),
    .X(_03263_));
 sky130_fd_sc_hd__o211a_1 _19300_ (.A1(\rbzero.spi_registers.new_texadd[3][17] ),
    .A2(_03254_),
    .B1(_03263_),
    .C1(_03252_),
    .X(_00872_));
 sky130_fd_sc_hd__or2_1 _19301_ (.A(\rbzero.spi_registers.texadd3[18] ),
    .B(_03255_),
    .X(_03264_));
 sky130_fd_sc_hd__buf_4 _19302_ (.A(_03212_),
    .X(_03265_));
 sky130_fd_sc_hd__o211a_1 _19303_ (.A1(\rbzero.spi_registers.new_texadd[3][18] ),
    .A2(_03254_),
    .B1(_03264_),
    .C1(_03265_),
    .X(_00873_));
 sky130_fd_sc_hd__or2_1 _19304_ (.A(\rbzero.spi_registers.texadd3[19] ),
    .B(_03255_),
    .X(_03266_));
 sky130_fd_sc_hd__o211a_1 _19305_ (.A1(\rbzero.spi_registers.new_texadd[3][19] ),
    .A2(_03254_),
    .B1(_03266_),
    .C1(_03265_),
    .X(_00874_));
 sky130_fd_sc_hd__or2_1 _19306_ (.A(\rbzero.spi_registers.texadd3[20] ),
    .B(_03241_),
    .X(_03267_));
 sky130_fd_sc_hd__o211a_1 _19307_ (.A1(\rbzero.spi_registers.new_texadd[3][20] ),
    .A2(_03239_),
    .B1(_03267_),
    .C1(_03265_),
    .X(_00875_));
 sky130_fd_sc_hd__or2_1 _19308_ (.A(\rbzero.spi_registers.texadd3[21] ),
    .B(_03241_),
    .X(_03268_));
 sky130_fd_sc_hd__o211a_1 _19309_ (.A1(\rbzero.spi_registers.new_texadd[3][21] ),
    .A2(_03239_),
    .B1(_03268_),
    .C1(_03265_),
    .X(_00876_));
 sky130_fd_sc_hd__or2_1 _19310_ (.A(\rbzero.spi_registers.texadd3[22] ),
    .B(_03241_),
    .X(_03269_));
 sky130_fd_sc_hd__o211a_1 _19311_ (.A1(\rbzero.spi_registers.new_texadd[3][22] ),
    .A2(_03239_),
    .B1(_03269_),
    .C1(_03265_),
    .X(_00877_));
 sky130_fd_sc_hd__or2_1 _19312_ (.A(\rbzero.spi_registers.texadd3[23] ),
    .B(_03241_),
    .X(_03270_));
 sky130_fd_sc_hd__o211a_1 _19313_ (.A1(\rbzero.spi_registers.new_texadd[3][23] ),
    .A2(_03239_),
    .B1(_03270_),
    .C1(_03265_),
    .X(_00878_));
 sky130_fd_sc_hd__nand2_2 _19314_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_03097_),
    .Y(_03271_));
 sky130_fd_sc_hd__and2_1 _19315_ (.A(\rbzero.spi_registers.got_new_leak ),
    .B(_03095_),
    .X(_03272_));
 sky130_fd_sc_hd__or2_1 _19316_ (.A(\rbzero.floor_leak[0] ),
    .B(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__o211a_1 _19317_ (.A1(\rbzero.spi_registers.new_leak[0] ),
    .A2(_03271_),
    .B1(_03273_),
    .C1(_03265_),
    .X(_00879_));
 sky130_fd_sc_hd__or2_1 _19318_ (.A(\rbzero.floor_leak[1] ),
    .B(_03272_),
    .X(_03274_));
 sky130_fd_sc_hd__o211a_1 _19319_ (.A1(\rbzero.spi_registers.new_leak[1] ),
    .A2(_03271_),
    .B1(_03274_),
    .C1(_03265_),
    .X(_00880_));
 sky130_fd_sc_hd__or2_1 _19320_ (.A(\rbzero.floor_leak[2] ),
    .B(_03272_),
    .X(_03275_));
 sky130_fd_sc_hd__o211a_1 _19321_ (.A1(\rbzero.spi_registers.new_leak[2] ),
    .A2(_03271_),
    .B1(_03275_),
    .C1(_03265_),
    .X(_00881_));
 sky130_fd_sc_hd__or2_1 _19322_ (.A(\rbzero.floor_leak[3] ),
    .B(_03272_),
    .X(_03276_));
 sky130_fd_sc_hd__o211a_1 _19323_ (.A1(\rbzero.spi_registers.new_leak[3] ),
    .A2(_03271_),
    .B1(_03276_),
    .C1(_03265_),
    .X(_00882_));
 sky130_fd_sc_hd__or2_1 _19324_ (.A(\rbzero.floor_leak[4] ),
    .B(_03272_),
    .X(_03277_));
 sky130_fd_sc_hd__clkbuf_4 _19325_ (.A(_03212_),
    .X(_03278_));
 sky130_fd_sc_hd__o211a_1 _19326_ (.A1(\rbzero.spi_registers.new_leak[4] ),
    .A2(_03271_),
    .B1(_03277_),
    .C1(_03278_),
    .X(_00883_));
 sky130_fd_sc_hd__or2_1 _19327_ (.A(\rbzero.floor_leak[5] ),
    .B(_03272_),
    .X(_03279_));
 sky130_fd_sc_hd__o211a_1 _19328_ (.A1(\rbzero.spi_registers.new_leak[5] ),
    .A2(_03271_),
    .B1(_03279_),
    .C1(_03278_),
    .X(_00884_));
 sky130_fd_sc_hd__nand2_2 _19329_ (.A(\rbzero.spi_registers.got_new_sky ),
    .B(_03097_),
    .Y(_03280_));
 sky130_fd_sc_hd__a31o_1 _19330_ (.A1(\rbzero.spi_registers.new_sky[0] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_03097_),
    .B1(_04409_),
    .X(_03281_));
 sky130_fd_sc_hd__a21o_1 _19331_ (.A1(\rbzero.color_sky[0] ),
    .A2(_03280_),
    .B1(_03281_),
    .X(_00885_));
 sky130_fd_sc_hd__and2_1 _19332_ (.A(\rbzero.spi_registers.got_new_sky ),
    .B(_03096_),
    .X(_03282_));
 sky130_fd_sc_hd__or2_1 _19333_ (.A(\rbzero.color_sky[1] ),
    .B(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__o211a_1 _19334_ (.A1(\rbzero.spi_registers.new_sky[1] ),
    .A2(_03280_),
    .B1(_03283_),
    .C1(_03278_),
    .X(_00886_));
 sky130_fd_sc_hd__a31o_1 _19335_ (.A1(\rbzero.spi_registers.new_sky[2] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_03097_),
    .B1(_04409_),
    .X(_03284_));
 sky130_fd_sc_hd__a21o_1 _19336_ (.A1(\rbzero.color_sky[2] ),
    .A2(_03280_),
    .B1(_03284_),
    .X(_00887_));
 sky130_fd_sc_hd__or2_1 _19337_ (.A(\rbzero.color_sky[3] ),
    .B(_03282_),
    .X(_03285_));
 sky130_fd_sc_hd__o211a_1 _19338_ (.A1(\rbzero.spi_registers.new_sky[3] ),
    .A2(_03280_),
    .B1(_03285_),
    .C1(_03278_),
    .X(_00888_));
 sky130_fd_sc_hd__a31o_1 _19339_ (.A1(\rbzero.spi_registers.new_sky[4] ),
    .A2(\rbzero.spi_registers.got_new_sky ),
    .A3(_03097_),
    .B1(_04409_),
    .X(_03286_));
 sky130_fd_sc_hd__a21o_1 _19340_ (.A1(\rbzero.color_sky[4] ),
    .A2(_03280_),
    .B1(_03286_),
    .X(_00889_));
 sky130_fd_sc_hd__or2_1 _19341_ (.A(\rbzero.color_sky[5] ),
    .B(_03282_),
    .X(_03287_));
 sky130_fd_sc_hd__o211a_1 _19342_ (.A1(\rbzero.spi_registers.new_sky[5] ),
    .A2(_03280_),
    .B1(_03287_),
    .C1(_03278_),
    .X(_00890_));
 sky130_fd_sc_hd__buf_4 _19343_ (.A(_03096_),
    .X(_03288_));
 sky130_fd_sc_hd__nand2_2 _19344_ (.A(\rbzero.spi_registers.got_new_floor ),
    .B(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__and2_1 _19345_ (.A(\rbzero.spi_registers.got_new_floor ),
    .B(_03096_),
    .X(_03290_));
 sky130_fd_sc_hd__or2_1 _19346_ (.A(\rbzero.color_floor[0] ),
    .B(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__o211a_1 _19347_ (.A1(\rbzero.spi_registers.new_floor[0] ),
    .A2(_03289_),
    .B1(_03291_),
    .C1(_03278_),
    .X(_00891_));
 sky130_fd_sc_hd__a31o_1 _19348_ (.A1(\rbzero.spi_registers.new_floor[1] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_03097_),
    .B1(_04409_),
    .X(_03292_));
 sky130_fd_sc_hd__a21o_1 _19349_ (.A1(\rbzero.color_floor[1] ),
    .A2(_03289_),
    .B1(_03292_),
    .X(_00892_));
 sky130_fd_sc_hd__or2_1 _19350_ (.A(\rbzero.color_floor[2] ),
    .B(_03290_),
    .X(_03293_));
 sky130_fd_sc_hd__o211a_1 _19351_ (.A1(\rbzero.spi_registers.new_floor[2] ),
    .A2(_03289_),
    .B1(_03293_),
    .C1(_03278_),
    .X(_00893_));
 sky130_fd_sc_hd__a31o_1 _19352_ (.A1(\rbzero.spi_registers.new_floor[3] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_03097_),
    .B1(_04409_),
    .X(_03294_));
 sky130_fd_sc_hd__a21o_1 _19353_ (.A1(\rbzero.color_floor[3] ),
    .A2(_03289_),
    .B1(_03294_),
    .X(_00894_));
 sky130_fd_sc_hd__or2_1 _19354_ (.A(\rbzero.color_floor[4] ),
    .B(_03290_),
    .X(_03295_));
 sky130_fd_sc_hd__o211a_1 _19355_ (.A1(\rbzero.spi_registers.new_floor[4] ),
    .A2(_03289_),
    .B1(_03295_),
    .C1(_03278_),
    .X(_00895_));
 sky130_fd_sc_hd__a31o_1 _19356_ (.A1(\rbzero.spi_registers.new_floor[5] ),
    .A2(\rbzero.spi_registers.got_new_floor ),
    .A3(_03097_),
    .B1(_04409_),
    .X(_03296_));
 sky130_fd_sc_hd__a21o_1 _19357_ (.A1(\rbzero.color_floor[5] ),
    .A2(_03289_),
    .B1(_03296_),
    .X(_00896_));
 sky130_fd_sc_hd__nand2_2 _19358_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_03097_),
    .Y(_03297_));
 sky130_fd_sc_hd__and2_1 _19359_ (.A(\rbzero.spi_registers.got_new_vshift ),
    .B(_03095_),
    .X(_03298_));
 sky130_fd_sc_hd__or2_1 _19360_ (.A(\rbzero.spi_registers.vshift[0] ),
    .B(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__o211a_1 _19361_ (.A1(\rbzero.spi_registers.new_vshift[0] ),
    .A2(_03297_),
    .B1(_03299_),
    .C1(_03278_),
    .X(_00897_));
 sky130_fd_sc_hd__or2_1 _19362_ (.A(\rbzero.spi_registers.vshift[1] ),
    .B(_03298_),
    .X(_03300_));
 sky130_fd_sc_hd__o211a_1 _19363_ (.A1(\rbzero.spi_registers.new_vshift[1] ),
    .A2(_03297_),
    .B1(_03300_),
    .C1(_03278_),
    .X(_00898_));
 sky130_fd_sc_hd__or2_1 _19364_ (.A(\rbzero.spi_registers.vshift[2] ),
    .B(_03298_),
    .X(_03301_));
 sky130_fd_sc_hd__buf_4 _19365_ (.A(_03212_),
    .X(_03302_));
 sky130_fd_sc_hd__o211a_1 _19366_ (.A1(\rbzero.spi_registers.new_vshift[2] ),
    .A2(_03297_),
    .B1(_03301_),
    .C1(_03302_),
    .X(_00899_));
 sky130_fd_sc_hd__or2_1 _19367_ (.A(\rbzero.spi_registers.vshift[3] ),
    .B(_03298_),
    .X(_03303_));
 sky130_fd_sc_hd__o211a_1 _19368_ (.A1(\rbzero.spi_registers.new_vshift[3] ),
    .A2(_03297_),
    .B1(_03303_),
    .C1(_03302_),
    .X(_00900_));
 sky130_fd_sc_hd__or2_1 _19369_ (.A(\rbzero.spi_registers.vshift[4] ),
    .B(_03298_),
    .X(_03304_));
 sky130_fd_sc_hd__o211a_1 _19370_ (.A1(\rbzero.spi_registers.new_vshift[4] ),
    .A2(_03297_),
    .B1(_03304_),
    .C1(_03302_),
    .X(_00901_));
 sky130_fd_sc_hd__or2_1 _19371_ (.A(\rbzero.spi_registers.vshift[5] ),
    .B(_03298_),
    .X(_03305_));
 sky130_fd_sc_hd__o211a_1 _19372_ (.A1(\rbzero.spi_registers.new_vshift[5] ),
    .A2(_03297_),
    .B1(_03305_),
    .C1(_03302_),
    .X(_00902_));
 sky130_fd_sc_hd__and4b_1 _19373_ (.A_N(\rbzero.spi_registers.spi_done ),
    .B(_02951_),
    .C(_02929_),
    .D(_02950_),
    .X(_03306_));
 sky130_fd_sc_hd__clkbuf_1 _19374_ (.A(_03306_),
    .X(_00903_));
 sky130_fd_sc_hd__or3b_1 _19375_ (.A(_02475_),
    .B(\rbzero.spi_registers.spi_cmd[3] ),
    .C_N(\rbzero.spi_registers.spi_done ),
    .X(_03307_));
 sky130_fd_sc_hd__or3_2 _19376_ (.A(_04408_),
    .B(_02930_),
    .C(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__buf_2 _19377_ (.A(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__mux2_1 _19378_ (.A0(_02473_),
    .A1(\rbzero.spi_registers.new_sky[0] ),
    .S(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__clkbuf_1 _19379_ (.A(_03310_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _19380_ (.A0(_02481_),
    .A1(\rbzero.spi_registers.new_sky[1] ),
    .S(_03309_),
    .X(_03311_));
 sky130_fd_sc_hd__clkbuf_1 _19381_ (.A(_03311_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _19382_ (.A0(_02483_),
    .A1(\rbzero.spi_registers.new_sky[2] ),
    .S(_03309_),
    .X(_03312_));
 sky130_fd_sc_hd__clkbuf_1 _19383_ (.A(_03312_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _19384_ (.A0(_02485_),
    .A1(\rbzero.spi_registers.new_sky[3] ),
    .S(_03309_),
    .X(_03313_));
 sky130_fd_sc_hd__clkbuf_1 _19385_ (.A(_03313_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _19386_ (.A0(_02487_),
    .A1(\rbzero.spi_registers.new_sky[4] ),
    .S(_03309_),
    .X(_03314_));
 sky130_fd_sc_hd__clkbuf_1 _19387_ (.A(_03314_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _19388_ (.A0(_02489_),
    .A1(\rbzero.spi_registers.new_sky[5] ),
    .S(_03309_),
    .X(_03315_));
 sky130_fd_sc_hd__clkbuf_1 _19389_ (.A(_03315_),
    .X(_00909_));
 sky130_fd_sc_hd__buf_4 _19390_ (.A(_03116_),
    .X(_03316_));
 sky130_fd_sc_hd__inv_2 _19391_ (.A(_03309_),
    .Y(_03317_));
 sky130_fd_sc_hd__a31o_1 _19392_ (.A1(\rbzero.spi_registers.got_new_sky ),
    .A2(_03118_),
    .A3(_03316_),
    .B1(_03317_),
    .X(_00910_));
 sky130_fd_sc_hd__or4b_2 _19393_ (.A(_02474_),
    .B(_04052_),
    .C(_03307_),
    .D_N(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_03318_));
 sky130_fd_sc_hd__buf_2 _19394_ (.A(_03318_),
    .X(_03319_));
 sky130_fd_sc_hd__mux2_1 _19395_ (.A0(_02473_),
    .A1(\rbzero.spi_registers.new_floor[0] ),
    .S(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__clkbuf_1 _19396_ (.A(_03320_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _19397_ (.A0(_02481_),
    .A1(\rbzero.spi_registers.new_floor[1] ),
    .S(_03319_),
    .X(_03321_));
 sky130_fd_sc_hd__clkbuf_1 _19398_ (.A(_03321_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _19399_ (.A0(_02483_),
    .A1(\rbzero.spi_registers.new_floor[2] ),
    .S(_03319_),
    .X(_03322_));
 sky130_fd_sc_hd__clkbuf_1 _19400_ (.A(_03322_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _19401_ (.A0(_02485_),
    .A1(\rbzero.spi_registers.new_floor[3] ),
    .S(_03319_),
    .X(_03323_));
 sky130_fd_sc_hd__clkbuf_1 _19402_ (.A(_03323_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _19403_ (.A0(_02487_),
    .A1(\rbzero.spi_registers.new_floor[4] ),
    .S(_03319_),
    .X(_03324_));
 sky130_fd_sc_hd__clkbuf_1 _19404_ (.A(_03324_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _19405_ (.A0(_02489_),
    .A1(\rbzero.spi_registers.new_floor[5] ),
    .S(_03319_),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_1 _19406_ (.A(_03325_),
    .X(_00916_));
 sky130_fd_sc_hd__inv_2 _19407_ (.A(_03319_),
    .Y(_03326_));
 sky130_fd_sc_hd__a31o_1 _19408_ (.A1(\rbzero.spi_registers.got_new_floor ),
    .A2(_03118_),
    .A3(_03316_),
    .B1(_03326_),
    .X(_00917_));
 sky130_fd_sc_hd__or2b_1 _19409_ (.A(\rbzero.spi_registers.spi_cmd[0] ),
    .B_N(_02474_),
    .X(_03327_));
 sky130_fd_sc_hd__or3_2 _19410_ (.A(_04408_),
    .B(_03307_),
    .C(_03327_),
    .X(_03328_));
 sky130_fd_sc_hd__buf_2 _19411_ (.A(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__mux2_1 _19412_ (.A0(_02473_),
    .A1(\rbzero.spi_registers.new_leak[0] ),
    .S(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__clkbuf_1 _19413_ (.A(_03330_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _19414_ (.A0(_02481_),
    .A1(\rbzero.spi_registers.new_leak[1] ),
    .S(_03329_),
    .X(_03331_));
 sky130_fd_sc_hd__clkbuf_1 _19415_ (.A(_03331_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _19416_ (.A0(_02483_),
    .A1(\rbzero.spi_registers.new_leak[2] ),
    .S(_03329_),
    .X(_03332_));
 sky130_fd_sc_hd__clkbuf_1 _19417_ (.A(_03332_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _19418_ (.A0(_02485_),
    .A1(\rbzero.spi_registers.new_leak[3] ),
    .S(_03329_),
    .X(_03333_));
 sky130_fd_sc_hd__clkbuf_1 _19419_ (.A(_03333_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _19420_ (.A0(_02487_),
    .A1(\rbzero.spi_registers.new_leak[4] ),
    .S(_03329_),
    .X(_03334_));
 sky130_fd_sc_hd__clkbuf_1 _19421_ (.A(_03334_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _19422_ (.A0(_02489_),
    .A1(\rbzero.spi_registers.new_leak[5] ),
    .S(_03329_),
    .X(_03335_));
 sky130_fd_sc_hd__clkbuf_1 _19423_ (.A(_03335_),
    .X(_00923_));
 sky130_fd_sc_hd__inv_2 _19424_ (.A(_03329_),
    .Y(_03336_));
 sky130_fd_sc_hd__a31o_1 _19425_ (.A1(\rbzero.spi_registers.got_new_leak ),
    .A2(_03118_),
    .A3(_03316_),
    .B1(_03336_),
    .X(_00924_));
 sky130_fd_sc_hd__or3_1 _19426_ (.A(_04408_),
    .B(_02932_),
    .C(_03307_),
    .X(_03337_));
 sky130_fd_sc_hd__clkbuf_4 _19427_ (.A(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__mux2_1 _19428_ (.A0(_02473_),
    .A1(\rbzero.spi_registers.new_other[0] ),
    .S(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__clkbuf_1 _19429_ (.A(_03339_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _19430_ (.A0(_02481_),
    .A1(\rbzero.spi_registers.new_other[1] ),
    .S(_03338_),
    .X(_03340_));
 sky130_fd_sc_hd__clkbuf_1 _19431_ (.A(_03340_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _19432_ (.A0(_02483_),
    .A1(\rbzero.spi_registers.new_other[2] ),
    .S(_03338_),
    .X(_03341_));
 sky130_fd_sc_hd__clkbuf_1 _19433_ (.A(_03341_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _19434_ (.A0(_02485_),
    .A1(\rbzero.spi_registers.new_other[3] ),
    .S(_03338_),
    .X(_03342_));
 sky130_fd_sc_hd__clkbuf_1 _19435_ (.A(_03342_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _19436_ (.A0(_02487_),
    .A1(\rbzero.spi_registers.new_other[4] ),
    .S(_03338_),
    .X(_03343_));
 sky130_fd_sc_hd__clkbuf_1 _19437_ (.A(_03343_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _19438_ (.A0(\rbzero.spi_registers.spi_buffer[6] ),
    .A1(\rbzero.spi_registers.new_other[6] ),
    .S(_03338_),
    .X(_03344_));
 sky130_fd_sc_hd__clkbuf_1 _19439_ (.A(_03344_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _19440_ (.A0(\rbzero.spi_registers.spi_buffer[7] ),
    .A1(\rbzero.spi_registers.new_other[7] ),
    .S(_03338_),
    .X(_03345_));
 sky130_fd_sc_hd__clkbuf_1 _19441_ (.A(_03345_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _19442_ (.A0(\rbzero.spi_registers.spi_buffer[8] ),
    .A1(\rbzero.spi_registers.new_other[8] ),
    .S(_03338_),
    .X(_03346_));
 sky130_fd_sc_hd__clkbuf_1 _19443_ (.A(_03346_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _19444_ (.A0(\rbzero.spi_registers.spi_buffer[9] ),
    .A1(\rbzero.spi_registers.new_other[9] ),
    .S(_03338_),
    .X(_03347_));
 sky130_fd_sc_hd__clkbuf_1 _19445_ (.A(_03347_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _19446_ (.A0(\rbzero.spi_registers.spi_buffer[10] ),
    .A1(\rbzero.spi_registers.new_other[10] ),
    .S(_03337_),
    .X(_03348_));
 sky130_fd_sc_hd__clkbuf_1 _19447_ (.A(_03348_),
    .X(_00934_));
 sky130_fd_sc_hd__inv_2 _19448_ (.A(_03338_),
    .Y(_03349_));
 sky130_fd_sc_hd__a31o_1 _19449_ (.A1(\rbzero.spi_registers.got_new_other ),
    .A2(_03118_),
    .A3(_03316_),
    .B1(_03349_),
    .X(_00935_));
 sky130_fd_sc_hd__and3_1 _19450_ (.A(\rbzero.spi_registers.spi_done ),
    .B(_02475_),
    .C(_02476_),
    .X(_03350_));
 sky130_fd_sc_hd__nor3b_4 _19451_ (.A(_04408_),
    .B(_02930_),
    .C_N(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__mux2_1 _19452_ (.A0(\rbzero.spi_registers.new_vshift[0] ),
    .A1(_02473_),
    .S(_03351_),
    .X(_03352_));
 sky130_fd_sc_hd__clkbuf_1 _19453_ (.A(_03352_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _19454_ (.A0(\rbzero.spi_registers.new_vshift[1] ),
    .A1(_02481_),
    .S(_03351_),
    .X(_03353_));
 sky130_fd_sc_hd__clkbuf_1 _19455_ (.A(_03353_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _19456_ (.A0(\rbzero.spi_registers.new_vshift[2] ),
    .A1(_02483_),
    .S(_03351_),
    .X(_03354_));
 sky130_fd_sc_hd__clkbuf_1 _19457_ (.A(_03354_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _19458_ (.A0(\rbzero.spi_registers.new_vshift[3] ),
    .A1(_02485_),
    .S(_03351_),
    .X(_03355_));
 sky130_fd_sc_hd__clkbuf_1 _19459_ (.A(_03355_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _19460_ (.A0(\rbzero.spi_registers.new_vshift[4] ),
    .A1(_02487_),
    .S(_03351_),
    .X(_03356_));
 sky130_fd_sc_hd__clkbuf_1 _19461_ (.A(_03356_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _19462_ (.A0(\rbzero.spi_registers.new_vshift[5] ),
    .A1(_02489_),
    .S(_03351_),
    .X(_03357_));
 sky130_fd_sc_hd__clkbuf_1 _19463_ (.A(_03357_),
    .X(_00941_));
 sky130_fd_sc_hd__a31o_1 _19464_ (.A1(\rbzero.spi_registers.got_new_vshift ),
    .A2(_03118_),
    .A3(_03316_),
    .B1(_03351_),
    .X(_00942_));
 sky130_fd_sc_hd__and4b_1 _19465_ (.A_N(_02474_),
    .B(_08116_),
    .C(_03350_),
    .D(\rbzero.spi_registers.spi_cmd[0] ),
    .X(_03358_));
 sky130_fd_sc_hd__mux2_1 _19466_ (.A0(\rbzero.spi_registers.new_vinf ),
    .A1(_02473_),
    .S(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__clkbuf_1 _19467_ (.A(_03359_),
    .X(_00943_));
 sky130_fd_sc_hd__a31o_1 _19468_ (.A1(\rbzero.spi_registers.got_new_vinf ),
    .A2(_03118_),
    .A3(_03316_),
    .B1(_03358_),
    .X(_00944_));
 sky130_fd_sc_hd__and4b_1 _19469_ (.A_N(\rbzero.spi_registers.spi_cmd[0] ),
    .B(_02474_),
    .C(_03974_),
    .D(_03350_),
    .X(_03360_));
 sky130_fd_sc_hd__clkbuf_4 _19470_ (.A(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__clkbuf_4 _19471_ (.A(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__mux2_1 _19472_ (.A0(\rbzero.spi_registers.new_mapd[0] ),
    .A1(_02473_),
    .S(_03362_),
    .X(_03363_));
 sky130_fd_sc_hd__clkbuf_1 _19473_ (.A(_03363_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _19474_ (.A0(\rbzero.spi_registers.new_mapd[1] ),
    .A1(_02481_),
    .S(_03362_),
    .X(_03364_));
 sky130_fd_sc_hd__clkbuf_1 _19475_ (.A(_03364_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _19476_ (.A0(\rbzero.spi_registers.new_mapd[2] ),
    .A1(_02483_),
    .S(_03362_),
    .X(_03365_));
 sky130_fd_sc_hd__clkbuf_1 _19477_ (.A(_03365_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _19478_ (.A0(\rbzero.spi_registers.new_mapd[3] ),
    .A1(_02485_),
    .S(_03362_),
    .X(_03366_));
 sky130_fd_sc_hd__clkbuf_1 _19479_ (.A(_03366_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _19480_ (.A0(\rbzero.spi_registers.new_mapd[4] ),
    .A1(_02487_),
    .S(_03362_),
    .X(_03367_));
 sky130_fd_sc_hd__clkbuf_1 _19481_ (.A(_03367_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _19482_ (.A0(\rbzero.spi_registers.new_mapd[5] ),
    .A1(_02489_),
    .S(_03362_),
    .X(_03368_));
 sky130_fd_sc_hd__clkbuf_1 _19483_ (.A(_03368_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _19484_ (.A0(\rbzero.spi_registers.new_mapd[6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03362_),
    .X(_03369_));
 sky130_fd_sc_hd__clkbuf_1 _19485_ (.A(_03369_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _19486_ (.A0(\rbzero.spi_registers.new_mapd[7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03362_),
    .X(_03370_));
 sky130_fd_sc_hd__clkbuf_1 _19487_ (.A(_03370_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _19488_ (.A0(\rbzero.spi_registers.new_mapd[8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03362_),
    .X(_03371_));
 sky130_fd_sc_hd__clkbuf_1 _19489_ (.A(_03371_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _19490_ (.A0(\rbzero.spi_registers.new_mapd[9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03361_),
    .X(_03372_));
 sky130_fd_sc_hd__clkbuf_1 _19491_ (.A(_03372_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _19492_ (.A0(\rbzero.spi_registers.new_mapd[10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03361_),
    .X(_03373_));
 sky130_fd_sc_hd__clkbuf_1 _19493_ (.A(_03373_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _19494_ (.A0(\rbzero.spi_registers.new_mapd[11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03361_),
    .X(_03374_));
 sky130_fd_sc_hd__clkbuf_1 _19495_ (.A(_03374_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _19496_ (.A0(\rbzero.spi_registers.new_mapd[12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03361_),
    .X(_03375_));
 sky130_fd_sc_hd__clkbuf_1 _19497_ (.A(_03375_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _19498_ (.A0(\rbzero.spi_registers.new_mapd[13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03361_),
    .X(_03376_));
 sky130_fd_sc_hd__clkbuf_1 _19499_ (.A(_03376_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _19500_ (.A0(\rbzero.spi_registers.new_mapd[14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03361_),
    .X(_03377_));
 sky130_fd_sc_hd__clkbuf_1 _19501_ (.A(_03377_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _19502_ (.A0(\rbzero.spi_registers.new_mapd[15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03361_),
    .X(_03378_));
 sky130_fd_sc_hd__clkbuf_1 _19503_ (.A(_03378_),
    .X(_00960_));
 sky130_fd_sc_hd__a31o_1 _19504_ (.A1(\rbzero.spi_registers.got_new_mapd ),
    .A2(_03118_),
    .A3(_03316_),
    .B1(_03362_),
    .X(_00961_));
 sky130_fd_sc_hd__and3_1 _19505_ (.A(_08116_),
    .B(_02936_),
    .C(_03350_),
    .X(_03379_));
 sky130_fd_sc_hd__clkbuf_4 _19506_ (.A(_03379_),
    .X(_03380_));
 sky130_fd_sc_hd__buf_4 _19507_ (.A(_03380_),
    .X(_03381_));
 sky130_fd_sc_hd__a31o_1 _19508_ (.A1(\rbzero.spi_registers.got_new_texadd[0] ),
    .A2(_08117_),
    .A3(_03316_),
    .B1(_03381_),
    .X(_00962_));
 sky130_fd_sc_hd__nor2_4 _19509_ (.A(_02477_),
    .B(_02930_),
    .Y(_03382_));
 sky130_fd_sc_hd__buf_4 _19510_ (.A(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__a31o_1 _19511_ (.A1(\rbzero.spi_registers.got_new_texadd[1] ),
    .A2(_08117_),
    .A3(_03316_),
    .B1(_03383_),
    .X(_00963_));
 sky130_fd_sc_hd__a31o_1 _19512_ (.A1(\rbzero.spi_registers.got_new_texadd[2] ),
    .A2(_08117_),
    .A3(_03316_),
    .B1(_02479_),
    .X(_00964_));
 sky130_fd_sc_hd__nor2_4 _19513_ (.A(_02477_),
    .B(_03327_),
    .Y(_03384_));
 sky130_fd_sc_hd__buf_4 _19514_ (.A(_03384_),
    .X(_03385_));
 sky130_fd_sc_hd__a31o_1 _19515_ (.A1(\rbzero.spi_registers.got_new_texadd[3] ),
    .A2(_08117_),
    .A3(_03116_),
    .B1(_03385_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _19516_ (.A0(\rbzero.spi_registers.new_texadd[0][0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_03381_),
    .X(_03386_));
 sky130_fd_sc_hd__clkbuf_1 _19517_ (.A(_03386_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _19518_ (.A0(\rbzero.spi_registers.new_texadd[0][1] ),
    .A1(_02481_),
    .S(_03381_),
    .X(_03387_));
 sky130_fd_sc_hd__clkbuf_1 _19519_ (.A(_03387_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _19520_ (.A0(\rbzero.spi_registers.new_texadd[0][2] ),
    .A1(_02483_),
    .S(_03381_),
    .X(_03388_));
 sky130_fd_sc_hd__clkbuf_1 _19521_ (.A(_03388_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _19522_ (.A0(\rbzero.spi_registers.new_texadd[0][3] ),
    .A1(_02485_),
    .S(_03381_),
    .X(_03389_));
 sky130_fd_sc_hd__clkbuf_1 _19523_ (.A(_03389_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _19524_ (.A0(\rbzero.spi_registers.new_texadd[0][4] ),
    .A1(_02487_),
    .S(_03381_),
    .X(_03390_));
 sky130_fd_sc_hd__clkbuf_1 _19525_ (.A(_03390_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _19526_ (.A0(\rbzero.spi_registers.new_texadd[0][5] ),
    .A1(_02489_),
    .S(_03381_),
    .X(_03391_));
 sky130_fd_sc_hd__clkbuf_1 _19527_ (.A(_03391_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _19528_ (.A0(\rbzero.spi_registers.new_texadd[0][6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03381_),
    .X(_03392_));
 sky130_fd_sc_hd__clkbuf_1 _19529_ (.A(_03392_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _19530_ (.A0(\rbzero.spi_registers.new_texadd[0][7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03381_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_1 _19531_ (.A(_03393_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _19532_ (.A0(\rbzero.spi_registers.new_texadd[0][8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03381_),
    .X(_03394_));
 sky130_fd_sc_hd__clkbuf_1 _19533_ (.A(_03394_),
    .X(_00974_));
 sky130_fd_sc_hd__buf_4 _19534_ (.A(_03380_),
    .X(_03395_));
 sky130_fd_sc_hd__mux2_1 _19535_ (.A0(\rbzero.spi_registers.new_texadd[0][9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03395_),
    .X(_03396_));
 sky130_fd_sc_hd__clkbuf_1 _19536_ (.A(_03396_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _19537_ (.A0(\rbzero.spi_registers.new_texadd[0][10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03395_),
    .X(_03397_));
 sky130_fd_sc_hd__clkbuf_1 _19538_ (.A(_03397_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _19539_ (.A0(\rbzero.spi_registers.new_texadd[0][11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03395_),
    .X(_03398_));
 sky130_fd_sc_hd__clkbuf_1 _19540_ (.A(_03398_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _19541_ (.A0(\rbzero.spi_registers.new_texadd[0][12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03395_),
    .X(_03399_));
 sky130_fd_sc_hd__clkbuf_1 _19542_ (.A(_03399_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _19543_ (.A0(\rbzero.spi_registers.new_texadd[0][13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03395_),
    .X(_03400_));
 sky130_fd_sc_hd__clkbuf_1 _19544_ (.A(_03400_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _19545_ (.A0(\rbzero.spi_registers.new_texadd[0][14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03395_),
    .X(_03401_));
 sky130_fd_sc_hd__clkbuf_1 _19546_ (.A(_03401_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _19547_ (.A0(\rbzero.spi_registers.new_texadd[0][15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03395_),
    .X(_03402_));
 sky130_fd_sc_hd__clkbuf_1 _19548_ (.A(_03402_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _19549_ (.A0(\rbzero.spi_registers.new_texadd[0][16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03395_),
    .X(_03403_));
 sky130_fd_sc_hd__clkbuf_1 _19550_ (.A(_03403_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _19551_ (.A0(\rbzero.spi_registers.new_texadd[0][17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03395_),
    .X(_03404_));
 sky130_fd_sc_hd__clkbuf_1 _19552_ (.A(_03404_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _19553_ (.A0(\rbzero.spi_registers.new_texadd[0][18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03395_),
    .X(_03405_));
 sky130_fd_sc_hd__clkbuf_1 _19554_ (.A(_03405_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _19555_ (.A0(\rbzero.spi_registers.new_texadd[0][19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03380_),
    .X(_03406_));
 sky130_fd_sc_hd__clkbuf_1 _19556_ (.A(_03406_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _19557_ (.A0(\rbzero.spi_registers.new_texadd[0][20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03380_),
    .X(_03407_));
 sky130_fd_sc_hd__clkbuf_1 _19558_ (.A(_03407_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _19559_ (.A0(\rbzero.spi_registers.new_texadd[0][21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03380_),
    .X(_03408_));
 sky130_fd_sc_hd__clkbuf_1 _19560_ (.A(_03408_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _19561_ (.A0(\rbzero.spi_registers.new_texadd[0][22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03380_),
    .X(_03409_));
 sky130_fd_sc_hd__clkbuf_1 _19562_ (.A(_03409_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _19563_ (.A0(\rbzero.spi_registers.new_texadd[0][23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_03380_),
    .X(_03410_));
 sky130_fd_sc_hd__clkbuf_1 _19564_ (.A(_03410_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _19565_ (.A0(\rbzero.spi_registers.new_texadd[1][0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_03383_),
    .X(_03411_));
 sky130_fd_sc_hd__clkbuf_1 _19566_ (.A(_03411_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _19567_ (.A0(\rbzero.spi_registers.new_texadd[1][1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_03383_),
    .X(_03412_));
 sky130_fd_sc_hd__clkbuf_1 _19568_ (.A(_03412_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _19569_ (.A0(\rbzero.spi_registers.new_texadd[1][2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_03383_),
    .X(_03413_));
 sky130_fd_sc_hd__clkbuf_1 _19570_ (.A(_03413_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _19571_ (.A0(\rbzero.spi_registers.new_texadd[1][3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_03383_),
    .X(_03414_));
 sky130_fd_sc_hd__clkbuf_1 _19572_ (.A(_03414_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _19573_ (.A0(\rbzero.spi_registers.new_texadd[1][4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_03383_),
    .X(_03415_));
 sky130_fd_sc_hd__clkbuf_1 _19574_ (.A(_03415_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _19575_ (.A0(\rbzero.spi_registers.new_texadd[1][5] ),
    .A1(_02489_),
    .S(_03383_),
    .X(_03416_));
 sky130_fd_sc_hd__clkbuf_1 _19576_ (.A(_03416_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _19577_ (.A0(\rbzero.spi_registers.new_texadd[1][6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03383_),
    .X(_03417_));
 sky130_fd_sc_hd__clkbuf_1 _19578_ (.A(_03417_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _19579_ (.A0(\rbzero.spi_registers.new_texadd[1][7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03383_),
    .X(_03418_));
 sky130_fd_sc_hd__clkbuf_1 _19580_ (.A(_03418_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _19581_ (.A0(\rbzero.spi_registers.new_texadd[1][8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03383_),
    .X(_03419_));
 sky130_fd_sc_hd__clkbuf_1 _19582_ (.A(_03419_),
    .X(_00998_));
 sky130_fd_sc_hd__buf_4 _19583_ (.A(_03382_),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_1 _19584_ (.A0(\rbzero.spi_registers.new_texadd[1][9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03420_),
    .X(_03421_));
 sky130_fd_sc_hd__clkbuf_1 _19585_ (.A(_03421_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _19586_ (.A0(\rbzero.spi_registers.new_texadd[1][10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03420_),
    .X(_03422_));
 sky130_fd_sc_hd__clkbuf_1 _19587_ (.A(_03422_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _19588_ (.A0(\rbzero.spi_registers.new_texadd[1][11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03420_),
    .X(_03423_));
 sky130_fd_sc_hd__clkbuf_1 _19589_ (.A(_03423_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _19590_ (.A0(\rbzero.spi_registers.new_texadd[1][12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03420_),
    .X(_03424_));
 sky130_fd_sc_hd__clkbuf_1 _19591_ (.A(_03424_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _19592_ (.A0(\rbzero.spi_registers.new_texadd[1][13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03420_),
    .X(_03425_));
 sky130_fd_sc_hd__clkbuf_1 _19593_ (.A(_03425_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _19594_ (.A0(\rbzero.spi_registers.new_texadd[1][14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03420_),
    .X(_03426_));
 sky130_fd_sc_hd__clkbuf_1 _19595_ (.A(_03426_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _19596_ (.A0(\rbzero.spi_registers.new_texadd[1][15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03420_),
    .X(_03427_));
 sky130_fd_sc_hd__clkbuf_1 _19597_ (.A(_03427_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _19598_ (.A0(\rbzero.spi_registers.new_texadd[1][16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03420_),
    .X(_03428_));
 sky130_fd_sc_hd__clkbuf_1 _19599_ (.A(_03428_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _19600_ (.A0(\rbzero.spi_registers.new_texadd[1][17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03420_),
    .X(_03429_));
 sky130_fd_sc_hd__clkbuf_1 _19601_ (.A(_03429_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _19602_ (.A0(\rbzero.spi_registers.new_texadd[1][18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03420_),
    .X(_03430_));
 sky130_fd_sc_hd__clkbuf_1 _19603_ (.A(_03430_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _19604_ (.A0(\rbzero.spi_registers.new_texadd[1][19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03382_),
    .X(_03431_));
 sky130_fd_sc_hd__clkbuf_1 _19605_ (.A(_03431_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _19606_ (.A0(\rbzero.spi_registers.new_texadd[1][20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03382_),
    .X(_03432_));
 sky130_fd_sc_hd__clkbuf_1 _19607_ (.A(_03432_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _19608_ (.A0(\rbzero.spi_registers.new_texadd[1][21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03382_),
    .X(_03433_));
 sky130_fd_sc_hd__clkbuf_1 _19609_ (.A(_03433_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _19610_ (.A0(\rbzero.spi_registers.new_texadd[1][22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03382_),
    .X(_03434_));
 sky130_fd_sc_hd__clkbuf_1 _19611_ (.A(_03434_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _19612_ (.A0(\rbzero.spi_registers.new_texadd[1][23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_03382_),
    .X(_03435_));
 sky130_fd_sc_hd__clkbuf_1 _19613_ (.A(_03435_),
    .X(_01013_));
 sky130_fd_sc_hd__or2_2 _19614_ (.A(net41),
    .B(net40),
    .X(_03436_));
 sky130_fd_sc_hd__nand2_1 _19615_ (.A(_03100_),
    .B(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__clkbuf_4 _19616_ (.A(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__o211a_1 _19617_ (.A1(\rbzero.pov.spi_done ),
    .A2(\rbzero.pov.ready ),
    .B1(_03118_),
    .C1(_03438_),
    .X(_01014_));
 sky130_fd_sc_hd__nor2b_2 _19618_ (.A(\rbzero.pov.sclk_buffer[2] ),
    .B_N(\rbzero.pov.sclk_buffer[1] ),
    .Y(_03439_));
 sky130_fd_sc_hd__nor2_2 _19619_ (.A(\rbzero.pov.ss_buffer[1] ),
    .B(_04052_),
    .Y(_03440_));
 sky130_fd_sc_hd__o21ai_1 _19620_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03439_),
    .B1(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__a21oi_1 _19621_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03439_),
    .B1(_03441_),
    .Y(_01015_));
 sky130_fd_sc_hd__and3_1 _19622_ (.A(\rbzero.pov.spi_counter[1] ),
    .B(\rbzero.pov.spi_counter[0] ),
    .C(_03439_),
    .X(_03442_));
 sky130_fd_sc_hd__a21o_1 _19623_ (.A1(\rbzero.pov.spi_counter[0] ),
    .A2(_03439_),
    .B1(\rbzero.pov.spi_counter[1] ),
    .X(_03443_));
 sky130_fd_sc_hd__and4bb_1 _19624_ (.A_N(\rbzero.pov.spi_counter[5] ),
    .B_N(\rbzero.pov.spi_counter[4] ),
    .C(\rbzero.pov.spi_counter[3] ),
    .D(\rbzero.pov.spi_counter[6] ),
    .X(_03444_));
 sky130_fd_sc_hd__and4bb_1 _19625_ (.A_N(\rbzero.pov.spi_counter[2] ),
    .B_N(\rbzero.pov.spi_counter[1] ),
    .C(\rbzero.pov.spi_counter[0] ),
    .D(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__a21boi_1 _19626_ (.A1(_03439_),
    .A2(_03445_),
    .B1_N(_03440_),
    .Y(_03446_));
 sky130_fd_sc_hd__and3b_1 _19627_ (.A_N(_03442_),
    .B(_03443_),
    .C(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_1 _19628_ (.A(_03447_),
    .X(_01016_));
 sky130_fd_sc_hd__and2_1 _19629_ (.A(\rbzero.pov.spi_counter[2] ),
    .B(_03442_),
    .X(_03448_));
 sky130_fd_sc_hd__o21ai_1 _19630_ (.A1(\rbzero.pov.spi_counter[2] ),
    .A2(_03442_),
    .B1(_03440_),
    .Y(_03449_));
 sky130_fd_sc_hd__nor2_1 _19631_ (.A(_03448_),
    .B(_03449_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _19632_ (.A(\rbzero.pov.spi_counter[3] ),
    .B(_03448_),
    .Y(_03450_));
 sky130_fd_sc_hd__o211a_1 _19633_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(_03448_),
    .B1(_03450_),
    .C1(_03446_),
    .X(_01018_));
 sky130_fd_sc_hd__and3_1 _19634_ (.A(\rbzero.pov.spi_counter[4] ),
    .B(\rbzero.pov.spi_counter[3] ),
    .C(_03448_),
    .X(_03451_));
 sky130_fd_sc_hd__a31o_1 _19635_ (.A1(\rbzero.pov.spi_counter[3] ),
    .A2(\rbzero.pov.spi_counter[2] ),
    .A3(_03442_),
    .B1(\rbzero.pov.spi_counter[4] ),
    .X(_03452_));
 sky130_fd_sc_hd__and3b_1 _19636_ (.A_N(_03451_),
    .B(_03440_),
    .C(_03452_),
    .X(_03453_));
 sky130_fd_sc_hd__clkbuf_1 _19637_ (.A(_03453_),
    .X(_01019_));
 sky130_fd_sc_hd__and2_1 _19638_ (.A(\rbzero.pov.spi_counter[5] ),
    .B(_03451_),
    .X(_03454_));
 sky130_fd_sc_hd__o21ai_1 _19639_ (.A1(\rbzero.pov.spi_counter[5] ),
    .A2(_03451_),
    .B1(_03440_),
    .Y(_03455_));
 sky130_fd_sc_hd__nor2_1 _19640_ (.A(_03454_),
    .B(_03455_),
    .Y(_01020_));
 sky130_fd_sc_hd__a21boi_1 _19641_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_03454_),
    .B1_N(_03446_),
    .Y(_03456_));
 sky130_fd_sc_hd__o21a_1 _19642_ (.A1(\rbzero.pov.spi_counter[6] ),
    .A2(_03454_),
    .B1(_03456_),
    .X(_01021_));
 sky130_fd_sc_hd__buf_1 _19643_ (.A(clknet_1_0__leaf__04634_),
    .X(_03457_));
 sky130_fd_sc_hd__buf_1 _19644_ (.A(clknet_1_1__leaf__03457_),
    .X(_03458_));
 sky130_fd_sc_hd__inv_2 _19646__28 (.A(clknet_1_1__leaf__03458_),
    .Y(net152));
 sky130_fd_sc_hd__inv_2 _19647__29 (.A(clknet_1_1__leaf__03458_),
    .Y(net153));
 sky130_fd_sc_hd__inv_2 _19648__30 (.A(clknet_1_1__leaf__03458_),
    .Y(net154));
 sky130_fd_sc_hd__inv_2 _19649__31 (.A(clknet_1_0__leaf__03458_),
    .Y(net155));
 sky130_fd_sc_hd__inv_2 _19650__32 (.A(clknet_1_0__leaf__03458_),
    .Y(net156));
 sky130_fd_sc_hd__inv_2 _19651__33 (.A(clknet_1_0__leaf__03458_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _19652__34 (.A(clknet_1_0__leaf__03458_),
    .Y(net158));
 sky130_fd_sc_hd__inv_2 _19653__35 (.A(clknet_1_0__leaf__03458_),
    .Y(net159));
 sky130_fd_sc_hd__inv_2 _19654__36 (.A(clknet_1_0__leaf__03458_),
    .Y(net160));
 sky130_fd_sc_hd__inv_2 _19656__37 (.A(clknet_1_0__leaf__03459_),
    .Y(net161));
 sky130_fd_sc_hd__buf_1 _19655_ (.A(clknet_1_0__leaf__03457_),
    .X(_03459_));
 sky130_fd_sc_hd__inv_2 _19657__38 (.A(clknet_1_0__leaf__03459_),
    .Y(net162));
 sky130_fd_sc_hd__inv_2 _19658__39 (.A(clknet_1_0__leaf__03459_),
    .Y(net163));
 sky130_fd_sc_hd__inv_2 _19659__40 (.A(clknet_1_0__leaf__03459_),
    .Y(net164));
 sky130_fd_sc_hd__inv_2 _19660__41 (.A(clknet_1_0__leaf__03459_),
    .Y(net165));
 sky130_fd_sc_hd__inv_2 _19661__42 (.A(clknet_1_0__leaf__03459_),
    .Y(net166));
 sky130_fd_sc_hd__inv_2 _19662__43 (.A(clknet_1_1__leaf__03459_),
    .Y(net167));
 sky130_fd_sc_hd__inv_2 _19663__44 (.A(clknet_1_1__leaf__03459_),
    .Y(net168));
 sky130_fd_sc_hd__inv_2 _19664__45 (.A(clknet_1_1__leaf__03459_),
    .Y(net169));
 sky130_fd_sc_hd__inv_2 _19665__46 (.A(clknet_1_1__leaf__03459_),
    .Y(net170));
 sky130_fd_sc_hd__inv_2 _19667__47 (.A(clknet_1_0__leaf__03460_),
    .Y(net171));
 sky130_fd_sc_hd__buf_1 _19666_ (.A(clknet_1_1__leaf__03457_),
    .X(_03460_));
 sky130_fd_sc_hd__inv_2 _19668__48 (.A(clknet_1_0__leaf__03460_),
    .Y(net172));
 sky130_fd_sc_hd__inv_2 _19669__49 (.A(clknet_1_0__leaf__03460_),
    .Y(net173));
 sky130_fd_sc_hd__inv_2 _19670__50 (.A(clknet_1_0__leaf__03460_),
    .Y(net174));
 sky130_fd_sc_hd__inv_2 _19671__51 (.A(clknet_1_0__leaf__03460_),
    .Y(net175));
 sky130_fd_sc_hd__inv_2 _19672__52 (.A(clknet_1_1__leaf__03460_),
    .Y(net176));
 sky130_fd_sc_hd__inv_2 _19673__53 (.A(clknet_1_1__leaf__03460_),
    .Y(net177));
 sky130_fd_sc_hd__inv_2 _19674__54 (.A(clknet_1_1__leaf__03460_),
    .Y(net178));
 sky130_fd_sc_hd__inv_2 _19675__55 (.A(clknet_1_1__leaf__03460_),
    .Y(net179));
 sky130_fd_sc_hd__inv_2 _19676__56 (.A(clknet_1_1__leaf__03460_),
    .Y(net180));
 sky130_fd_sc_hd__inv_2 _19678__57 (.A(clknet_1_1__leaf__03461_),
    .Y(net181));
 sky130_fd_sc_hd__buf_1 _19677_ (.A(clknet_1_0__leaf__03457_),
    .X(_03461_));
 sky130_fd_sc_hd__inv_2 _19679__58 (.A(clknet_1_1__leaf__03461_),
    .Y(net182));
 sky130_fd_sc_hd__inv_2 _19680__59 (.A(clknet_1_1__leaf__03461_),
    .Y(net183));
 sky130_fd_sc_hd__inv_2 _19681__60 (.A(clknet_1_1__leaf__03461_),
    .Y(net184));
 sky130_fd_sc_hd__inv_2 _19682__61 (.A(clknet_1_1__leaf__03461_),
    .Y(net185));
 sky130_fd_sc_hd__inv_2 _19683__62 (.A(clknet_1_1__leaf__03461_),
    .Y(net186));
 sky130_fd_sc_hd__inv_2 _19684__63 (.A(clknet_1_0__leaf__03461_),
    .Y(net187));
 sky130_fd_sc_hd__inv_2 _19685__64 (.A(clknet_1_0__leaf__03461_),
    .Y(net188));
 sky130_fd_sc_hd__inv_2 _19686__65 (.A(clknet_1_0__leaf__03461_),
    .Y(net189));
 sky130_fd_sc_hd__inv_2 _19687__66 (.A(clknet_1_0__leaf__03461_),
    .Y(net190));
 sky130_fd_sc_hd__inv_2 _19689__67 (.A(clknet_1_1__leaf__03462_),
    .Y(net191));
 sky130_fd_sc_hd__buf_1 _19688_ (.A(clknet_1_0__leaf__03457_),
    .X(_03462_));
 sky130_fd_sc_hd__inv_2 _19690__68 (.A(clknet_1_1__leaf__03462_),
    .Y(net192));
 sky130_fd_sc_hd__inv_2 _19691__69 (.A(clknet_1_0__leaf__03462_),
    .Y(net193));
 sky130_fd_sc_hd__inv_2 _19692__70 (.A(clknet_1_0__leaf__03462_),
    .Y(net194));
 sky130_fd_sc_hd__inv_2 _19693__71 (.A(clknet_1_0__leaf__03462_),
    .Y(net195));
 sky130_fd_sc_hd__inv_2 _19694__72 (.A(clknet_1_0__leaf__03462_),
    .Y(net196));
 sky130_fd_sc_hd__inv_2 _19695__73 (.A(clknet_1_0__leaf__03462_),
    .Y(net197));
 sky130_fd_sc_hd__inv_2 _19696__74 (.A(clknet_1_1__leaf__03462_),
    .Y(net198));
 sky130_fd_sc_hd__inv_2 _19697__75 (.A(clknet_1_1__leaf__03462_),
    .Y(net199));
 sky130_fd_sc_hd__inv_2 _19698__76 (.A(clknet_1_1__leaf__03462_),
    .Y(net200));
 sky130_fd_sc_hd__inv_2 _19700__77 (.A(clknet_1_0__leaf__03463_),
    .Y(net201));
 sky130_fd_sc_hd__buf_1 _19699_ (.A(clknet_1_0__leaf__03457_),
    .X(_03463_));
 sky130_fd_sc_hd__inv_2 _19701__78 (.A(clknet_1_0__leaf__03463_),
    .Y(net202));
 sky130_fd_sc_hd__inv_2 _19702__79 (.A(clknet_1_0__leaf__03463_),
    .Y(net203));
 sky130_fd_sc_hd__inv_2 _19703__80 (.A(clknet_1_0__leaf__03463_),
    .Y(net204));
 sky130_fd_sc_hd__inv_2 _19704__81 (.A(clknet_1_0__leaf__03463_),
    .Y(net205));
 sky130_fd_sc_hd__inv_2 _19705__82 (.A(clknet_1_1__leaf__03463_),
    .Y(net206));
 sky130_fd_sc_hd__inv_2 _19706__83 (.A(clknet_1_1__leaf__03463_),
    .Y(net207));
 sky130_fd_sc_hd__inv_2 _19707__84 (.A(clknet_1_1__leaf__03463_),
    .Y(net208));
 sky130_fd_sc_hd__inv_2 _19708__85 (.A(clknet_1_1__leaf__03463_),
    .Y(net209));
 sky130_fd_sc_hd__inv_2 _19709__86 (.A(clknet_1_1__leaf__03463_),
    .Y(net210));
 sky130_fd_sc_hd__inv_2 _19712__87 (.A(clknet_1_0__leaf__03465_),
    .Y(net211));
 sky130_fd_sc_hd__buf_1 _19710_ (.A(clknet_1_1__leaf__04634_),
    .X(_03464_));
 sky130_fd_sc_hd__buf_1 _19711_ (.A(clknet_1_0__leaf__03464_),
    .X(_03465_));
 sky130_fd_sc_hd__inv_2 _19713__88 (.A(clknet_1_0__leaf__03465_),
    .Y(net212));
 sky130_fd_sc_hd__inv_2 _19714__89 (.A(clknet_1_0__leaf__03465_),
    .Y(net213));
 sky130_fd_sc_hd__inv_2 _19715__90 (.A(clknet_1_0__leaf__03465_),
    .Y(net214));
 sky130_fd_sc_hd__inv_2 _20218__91 (.A(clknet_1_1__leaf__03465_),
    .Y(net215));
 sky130_fd_sc_hd__nand2_1 _19716_ (.A(_03440_),
    .B(_03439_),
    .Y(_03466_));
 sky130_fd_sc_hd__clkbuf_4 _19717_ (.A(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__clkbuf_4 _19718_ (.A(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__mux2_1 _19719_ (.A0(\rbzero.pov.mosi ),
    .A1(\rbzero.pov.spi_buffer[0] ),
    .S(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__clkbuf_1 _19720_ (.A(_03469_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _19721_ (.A0(\rbzero.pov.spi_buffer[0] ),
    .A1(\rbzero.pov.spi_buffer[1] ),
    .S(_03468_),
    .X(_03470_));
 sky130_fd_sc_hd__clkbuf_1 _19722_ (.A(_03470_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _19723_ (.A0(\rbzero.pov.spi_buffer[1] ),
    .A1(\rbzero.pov.spi_buffer[2] ),
    .S(_03468_),
    .X(_03471_));
 sky130_fd_sc_hd__clkbuf_1 _19724_ (.A(_03471_),
    .X(_01088_));
 sky130_fd_sc_hd__mux2_1 _19725_ (.A0(\rbzero.pov.spi_buffer[2] ),
    .A1(\rbzero.pov.spi_buffer[3] ),
    .S(_03468_),
    .X(_03472_));
 sky130_fd_sc_hd__clkbuf_1 _19726_ (.A(_03472_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _19727_ (.A0(\rbzero.pov.spi_buffer[3] ),
    .A1(\rbzero.pov.spi_buffer[4] ),
    .S(_03468_),
    .X(_03473_));
 sky130_fd_sc_hd__clkbuf_1 _19728_ (.A(_03473_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _19729_ (.A0(\rbzero.pov.spi_buffer[4] ),
    .A1(\rbzero.pov.spi_buffer[5] ),
    .S(_03468_),
    .X(_03474_));
 sky130_fd_sc_hd__clkbuf_1 _19730_ (.A(_03474_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _19731_ (.A0(\rbzero.pov.spi_buffer[5] ),
    .A1(\rbzero.pov.spi_buffer[6] ),
    .S(_03468_),
    .X(_03475_));
 sky130_fd_sc_hd__clkbuf_1 _19732_ (.A(_03475_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _19733_ (.A0(net511),
    .A1(\rbzero.pov.spi_buffer[7] ),
    .S(_03468_),
    .X(_03476_));
 sky130_fd_sc_hd__clkbuf_1 _19734_ (.A(_03476_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _19735_ (.A0(\rbzero.pov.spi_buffer[7] ),
    .A1(\rbzero.pov.spi_buffer[8] ),
    .S(_03468_),
    .X(_03477_));
 sky130_fd_sc_hd__clkbuf_1 _19736_ (.A(_03477_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _19737_ (.A0(\rbzero.pov.spi_buffer[8] ),
    .A1(\rbzero.pov.spi_buffer[9] ),
    .S(_03468_),
    .X(_03478_));
 sky130_fd_sc_hd__clkbuf_1 _19738_ (.A(_03478_),
    .X(_01095_));
 sky130_fd_sc_hd__clkbuf_4 _19739_ (.A(_03467_),
    .X(_03479_));
 sky130_fd_sc_hd__mux2_1 _19740_ (.A0(\rbzero.pov.spi_buffer[9] ),
    .A1(\rbzero.pov.spi_buffer[10] ),
    .S(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__clkbuf_1 _19741_ (.A(_03480_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _19742_ (.A0(\rbzero.pov.spi_buffer[10] ),
    .A1(\rbzero.pov.spi_buffer[11] ),
    .S(_03479_),
    .X(_03481_));
 sky130_fd_sc_hd__clkbuf_1 _19743_ (.A(_03481_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _19744_ (.A0(\rbzero.pov.spi_buffer[11] ),
    .A1(\rbzero.pov.spi_buffer[12] ),
    .S(_03479_),
    .X(_03482_));
 sky130_fd_sc_hd__clkbuf_1 _19745_ (.A(_03482_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _19746_ (.A0(\rbzero.pov.spi_buffer[12] ),
    .A1(\rbzero.pov.spi_buffer[13] ),
    .S(_03479_),
    .X(_03483_));
 sky130_fd_sc_hd__clkbuf_1 _19747_ (.A(_03483_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _19748_ (.A0(\rbzero.pov.spi_buffer[13] ),
    .A1(\rbzero.pov.spi_buffer[14] ),
    .S(_03479_),
    .X(_03484_));
 sky130_fd_sc_hd__clkbuf_1 _19749_ (.A(_03484_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _19750_ (.A0(\rbzero.pov.spi_buffer[14] ),
    .A1(\rbzero.pov.spi_buffer[15] ),
    .S(_03479_),
    .X(_03485_));
 sky130_fd_sc_hd__clkbuf_1 _19751_ (.A(_03485_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _19752_ (.A0(\rbzero.pov.spi_buffer[15] ),
    .A1(\rbzero.pov.spi_buffer[16] ),
    .S(_03479_),
    .X(_03486_));
 sky130_fd_sc_hd__clkbuf_1 _19753_ (.A(_03486_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _19754_ (.A0(\rbzero.pov.spi_buffer[16] ),
    .A1(\rbzero.pov.spi_buffer[17] ),
    .S(_03479_),
    .X(_03487_));
 sky130_fd_sc_hd__clkbuf_1 _19755_ (.A(_03487_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _19756_ (.A0(\rbzero.pov.spi_buffer[17] ),
    .A1(\rbzero.pov.spi_buffer[18] ),
    .S(_03479_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_1 _19757_ (.A(_03488_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _19758_ (.A0(\rbzero.pov.spi_buffer[18] ),
    .A1(\rbzero.pov.spi_buffer[19] ),
    .S(_03479_),
    .X(_03489_));
 sky130_fd_sc_hd__clkbuf_1 _19759_ (.A(_03489_),
    .X(_01105_));
 sky130_fd_sc_hd__clkbuf_4 _19760_ (.A(_03467_),
    .X(_03490_));
 sky130_fd_sc_hd__mux2_1 _19761_ (.A0(\rbzero.pov.spi_buffer[19] ),
    .A1(\rbzero.pov.spi_buffer[20] ),
    .S(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__clkbuf_1 _19762_ (.A(_03491_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _19763_ (.A0(\rbzero.pov.spi_buffer[20] ),
    .A1(\rbzero.pov.spi_buffer[21] ),
    .S(_03490_),
    .X(_03492_));
 sky130_fd_sc_hd__clkbuf_1 _19764_ (.A(_03492_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _19765_ (.A0(\rbzero.pov.spi_buffer[21] ),
    .A1(\rbzero.pov.spi_buffer[22] ),
    .S(_03490_),
    .X(_03493_));
 sky130_fd_sc_hd__clkbuf_1 _19766_ (.A(_03493_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _19767_ (.A0(\rbzero.pov.spi_buffer[22] ),
    .A1(\rbzero.pov.spi_buffer[23] ),
    .S(_03490_),
    .X(_03494_));
 sky130_fd_sc_hd__clkbuf_1 _19768_ (.A(_03494_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _19769_ (.A0(\rbzero.pov.spi_buffer[23] ),
    .A1(\rbzero.pov.spi_buffer[24] ),
    .S(_03490_),
    .X(_03495_));
 sky130_fd_sc_hd__clkbuf_1 _19770_ (.A(_03495_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _19771_ (.A0(\rbzero.pov.spi_buffer[24] ),
    .A1(\rbzero.pov.spi_buffer[25] ),
    .S(_03490_),
    .X(_03496_));
 sky130_fd_sc_hd__clkbuf_1 _19772_ (.A(_03496_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _19773_ (.A0(\rbzero.pov.spi_buffer[25] ),
    .A1(\rbzero.pov.spi_buffer[26] ),
    .S(_03490_),
    .X(_03497_));
 sky130_fd_sc_hd__clkbuf_1 _19774_ (.A(_03497_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _19775_ (.A0(\rbzero.pov.spi_buffer[26] ),
    .A1(\rbzero.pov.spi_buffer[27] ),
    .S(_03490_),
    .X(_03498_));
 sky130_fd_sc_hd__clkbuf_1 _19776_ (.A(_03498_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _19777_ (.A0(\rbzero.pov.spi_buffer[27] ),
    .A1(\rbzero.pov.spi_buffer[28] ),
    .S(_03490_),
    .X(_03499_));
 sky130_fd_sc_hd__clkbuf_1 _19778_ (.A(_03499_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _19779_ (.A0(\rbzero.pov.spi_buffer[28] ),
    .A1(\rbzero.pov.spi_buffer[29] ),
    .S(_03490_),
    .X(_03500_));
 sky130_fd_sc_hd__clkbuf_1 _19780_ (.A(_03500_),
    .X(_01115_));
 sky130_fd_sc_hd__clkbuf_4 _19781_ (.A(_03467_),
    .X(_03501_));
 sky130_fd_sc_hd__mux2_1 _19782_ (.A0(\rbzero.pov.spi_buffer[29] ),
    .A1(\rbzero.pov.spi_buffer[30] ),
    .S(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__clkbuf_1 _19783_ (.A(_03502_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _19784_ (.A0(\rbzero.pov.spi_buffer[30] ),
    .A1(\rbzero.pov.spi_buffer[31] ),
    .S(_03501_),
    .X(_03503_));
 sky130_fd_sc_hd__clkbuf_1 _19785_ (.A(_03503_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _19786_ (.A0(\rbzero.pov.spi_buffer[31] ),
    .A1(\rbzero.pov.spi_buffer[32] ),
    .S(_03501_),
    .X(_03504_));
 sky130_fd_sc_hd__clkbuf_1 _19787_ (.A(_03504_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _19788_ (.A0(\rbzero.pov.spi_buffer[32] ),
    .A1(\rbzero.pov.spi_buffer[33] ),
    .S(_03501_),
    .X(_03505_));
 sky130_fd_sc_hd__clkbuf_1 _19789_ (.A(_03505_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _19790_ (.A0(\rbzero.pov.spi_buffer[33] ),
    .A1(\rbzero.pov.spi_buffer[34] ),
    .S(_03501_),
    .X(_03506_));
 sky130_fd_sc_hd__clkbuf_1 _19791_ (.A(_03506_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _19792_ (.A0(\rbzero.pov.spi_buffer[34] ),
    .A1(\rbzero.pov.spi_buffer[35] ),
    .S(_03501_),
    .X(_03507_));
 sky130_fd_sc_hd__clkbuf_1 _19793_ (.A(_03507_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _19794_ (.A0(\rbzero.pov.spi_buffer[35] ),
    .A1(\rbzero.pov.spi_buffer[36] ),
    .S(_03501_),
    .X(_03508_));
 sky130_fd_sc_hd__clkbuf_1 _19795_ (.A(_03508_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _19796_ (.A0(\rbzero.pov.spi_buffer[36] ),
    .A1(\rbzero.pov.spi_buffer[37] ),
    .S(_03501_),
    .X(_03509_));
 sky130_fd_sc_hd__clkbuf_1 _19797_ (.A(_03509_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _19798_ (.A0(\rbzero.pov.spi_buffer[37] ),
    .A1(\rbzero.pov.spi_buffer[38] ),
    .S(_03501_),
    .X(_03510_));
 sky130_fd_sc_hd__clkbuf_1 _19799_ (.A(_03510_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _19800_ (.A0(\rbzero.pov.spi_buffer[38] ),
    .A1(\rbzero.pov.spi_buffer[39] ),
    .S(_03501_),
    .X(_03511_));
 sky130_fd_sc_hd__clkbuf_1 _19801_ (.A(_03511_),
    .X(_01125_));
 sky130_fd_sc_hd__buf_4 _19802_ (.A(_03467_),
    .X(_03512_));
 sky130_fd_sc_hd__mux2_1 _19803_ (.A0(\rbzero.pov.spi_buffer[39] ),
    .A1(\rbzero.pov.spi_buffer[40] ),
    .S(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__clkbuf_1 _19804_ (.A(_03513_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _19805_ (.A0(\rbzero.pov.spi_buffer[40] ),
    .A1(\rbzero.pov.spi_buffer[41] ),
    .S(_03512_),
    .X(_03514_));
 sky130_fd_sc_hd__clkbuf_1 _19806_ (.A(_03514_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _19807_ (.A0(\rbzero.pov.spi_buffer[41] ),
    .A1(\rbzero.pov.spi_buffer[42] ),
    .S(_03512_),
    .X(_03515_));
 sky130_fd_sc_hd__clkbuf_1 _19808_ (.A(_03515_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _19809_ (.A0(\rbzero.pov.spi_buffer[42] ),
    .A1(\rbzero.pov.spi_buffer[43] ),
    .S(_03512_),
    .X(_03516_));
 sky130_fd_sc_hd__clkbuf_1 _19810_ (.A(_03516_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _19811_ (.A0(\rbzero.pov.spi_buffer[43] ),
    .A1(\rbzero.pov.spi_buffer[44] ),
    .S(_03512_),
    .X(_03517_));
 sky130_fd_sc_hd__clkbuf_1 _19812_ (.A(_03517_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _19813_ (.A0(\rbzero.pov.spi_buffer[44] ),
    .A1(\rbzero.pov.spi_buffer[45] ),
    .S(_03512_),
    .X(_03518_));
 sky130_fd_sc_hd__clkbuf_1 _19814_ (.A(_03518_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _19815_ (.A0(\rbzero.pov.spi_buffer[45] ),
    .A1(\rbzero.pov.spi_buffer[46] ),
    .S(_03512_),
    .X(_03519_));
 sky130_fd_sc_hd__clkbuf_1 _19816_ (.A(_03519_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _19817_ (.A0(\rbzero.pov.spi_buffer[46] ),
    .A1(\rbzero.pov.spi_buffer[47] ),
    .S(_03512_),
    .X(_03520_));
 sky130_fd_sc_hd__clkbuf_1 _19818_ (.A(_03520_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _19819_ (.A0(\rbzero.pov.spi_buffer[47] ),
    .A1(\rbzero.pov.spi_buffer[48] ),
    .S(_03512_),
    .X(_03521_));
 sky130_fd_sc_hd__clkbuf_1 _19820_ (.A(_03521_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _19821_ (.A0(\rbzero.pov.spi_buffer[48] ),
    .A1(\rbzero.pov.spi_buffer[49] ),
    .S(_03512_),
    .X(_03522_));
 sky130_fd_sc_hd__clkbuf_1 _19822_ (.A(_03522_),
    .X(_01135_));
 sky130_fd_sc_hd__clkbuf_4 _19823_ (.A(_03467_),
    .X(_03523_));
 sky130_fd_sc_hd__mux2_1 _19824_ (.A0(\rbzero.pov.spi_buffer[49] ),
    .A1(\rbzero.pov.spi_buffer[50] ),
    .S(_03523_),
    .X(_03524_));
 sky130_fd_sc_hd__clkbuf_1 _19825_ (.A(_03524_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _19826_ (.A0(\rbzero.pov.spi_buffer[50] ),
    .A1(\rbzero.pov.spi_buffer[51] ),
    .S(_03523_),
    .X(_03525_));
 sky130_fd_sc_hd__clkbuf_1 _19827_ (.A(_03525_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _19828_ (.A0(\rbzero.pov.spi_buffer[51] ),
    .A1(\rbzero.pov.spi_buffer[52] ),
    .S(_03523_),
    .X(_03526_));
 sky130_fd_sc_hd__clkbuf_1 _19829_ (.A(_03526_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _19830_ (.A0(\rbzero.pov.spi_buffer[52] ),
    .A1(\rbzero.pov.spi_buffer[53] ),
    .S(_03523_),
    .X(_03527_));
 sky130_fd_sc_hd__clkbuf_1 _19831_ (.A(_03527_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _19832_ (.A0(\rbzero.pov.spi_buffer[53] ),
    .A1(\rbzero.pov.spi_buffer[54] ),
    .S(_03523_),
    .X(_03528_));
 sky130_fd_sc_hd__clkbuf_1 _19833_ (.A(_03528_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _19834_ (.A0(\rbzero.pov.spi_buffer[54] ),
    .A1(\rbzero.pov.spi_buffer[55] ),
    .S(_03523_),
    .X(_03529_));
 sky130_fd_sc_hd__clkbuf_1 _19835_ (.A(_03529_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _19836_ (.A0(\rbzero.pov.spi_buffer[55] ),
    .A1(\rbzero.pov.spi_buffer[56] ),
    .S(_03523_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_1 _19837_ (.A(_03530_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _19838_ (.A0(\rbzero.pov.spi_buffer[56] ),
    .A1(\rbzero.pov.spi_buffer[57] ),
    .S(_03523_),
    .X(_03531_));
 sky130_fd_sc_hd__clkbuf_1 _19839_ (.A(_03531_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _19840_ (.A0(\rbzero.pov.spi_buffer[57] ),
    .A1(\rbzero.pov.spi_buffer[58] ),
    .S(_03523_),
    .X(_03532_));
 sky130_fd_sc_hd__clkbuf_1 _19841_ (.A(_03532_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _19842_ (.A0(\rbzero.pov.spi_buffer[58] ),
    .A1(\rbzero.pov.spi_buffer[59] ),
    .S(_03523_),
    .X(_03533_));
 sky130_fd_sc_hd__clkbuf_1 _19843_ (.A(_03533_),
    .X(_01145_));
 sky130_fd_sc_hd__buf_4 _19844_ (.A(_03466_),
    .X(_03534_));
 sky130_fd_sc_hd__mux2_1 _19845_ (.A0(\rbzero.pov.spi_buffer[59] ),
    .A1(\rbzero.pov.spi_buffer[60] ),
    .S(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__clkbuf_1 _19846_ (.A(_03535_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _19847_ (.A0(\rbzero.pov.spi_buffer[60] ),
    .A1(\rbzero.pov.spi_buffer[61] ),
    .S(_03534_),
    .X(_03536_));
 sky130_fd_sc_hd__clkbuf_1 _19848_ (.A(_03536_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _19849_ (.A0(\rbzero.pov.spi_buffer[61] ),
    .A1(\rbzero.pov.spi_buffer[62] ),
    .S(_03534_),
    .X(_03537_));
 sky130_fd_sc_hd__clkbuf_1 _19850_ (.A(_03537_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _19851_ (.A0(\rbzero.pov.spi_buffer[62] ),
    .A1(\rbzero.pov.spi_buffer[63] ),
    .S(_03534_),
    .X(_03538_));
 sky130_fd_sc_hd__clkbuf_1 _19852_ (.A(_03538_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _19853_ (.A0(\rbzero.pov.spi_buffer[63] ),
    .A1(\rbzero.pov.spi_buffer[64] ),
    .S(_03534_),
    .X(_03539_));
 sky130_fd_sc_hd__clkbuf_1 _19854_ (.A(_03539_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _19855_ (.A0(\rbzero.pov.spi_buffer[64] ),
    .A1(\rbzero.pov.spi_buffer[65] ),
    .S(_03534_),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_1 _19856_ (.A(_03540_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _19857_ (.A0(\rbzero.pov.spi_buffer[65] ),
    .A1(\rbzero.pov.spi_buffer[66] ),
    .S(_03534_),
    .X(_03541_));
 sky130_fd_sc_hd__clkbuf_1 _19858_ (.A(_03541_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _19859_ (.A0(\rbzero.pov.spi_buffer[66] ),
    .A1(\rbzero.pov.spi_buffer[67] ),
    .S(_03534_),
    .X(_03542_));
 sky130_fd_sc_hd__clkbuf_1 _19860_ (.A(_03542_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _19861_ (.A0(\rbzero.pov.spi_buffer[67] ),
    .A1(\rbzero.pov.spi_buffer[68] ),
    .S(_03534_),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_1 _19862_ (.A(_03543_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _19863_ (.A0(\rbzero.pov.spi_buffer[68] ),
    .A1(\rbzero.pov.spi_buffer[69] ),
    .S(_03534_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_1 _19864_ (.A(_03544_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _19865_ (.A0(\rbzero.pov.spi_buffer[69] ),
    .A1(\rbzero.pov.spi_buffer[70] ),
    .S(_03467_),
    .X(_03545_));
 sky130_fd_sc_hd__clkbuf_1 _19866_ (.A(_03545_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _19867_ (.A0(\rbzero.pov.spi_buffer[70] ),
    .A1(\rbzero.pov.spi_buffer[71] ),
    .S(_03467_),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_1 _19868_ (.A(_03546_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _19869_ (.A0(\rbzero.pov.spi_buffer[71] ),
    .A1(\rbzero.pov.spi_buffer[72] ),
    .S(_03467_),
    .X(_03547_));
 sky130_fd_sc_hd__clkbuf_1 _19870_ (.A(_03547_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _19871_ (.A0(\rbzero.pov.spi_buffer[72] ),
    .A1(\rbzero.pov.spi_buffer[73] ),
    .S(_03467_),
    .X(_03548_));
 sky130_fd_sc_hd__clkbuf_1 _19872_ (.A(_03548_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _19873_ (.A0(_05711_),
    .A1(\rbzero.pov.mosi_buffer[0] ),
    .S(_09734_),
    .X(_03549_));
 sky130_fd_sc_hd__clkbuf_1 _19874_ (.A(_03549_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _19875_ (.A0(\rbzero.pov.mosi ),
    .A1(\rbzero.pov.mosi_buffer[0] ),
    .S(_03084_),
    .X(_03550_));
 sky130_fd_sc_hd__clkbuf_1 _19876_ (.A(_03550_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _19877_ (.A0(net53),
    .A1(\rbzero.pov.ss_buffer[0] ),
    .S(_09734_),
    .X(_03551_));
 sky130_fd_sc_hd__clkbuf_1 _19878_ (.A(_03551_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _19879_ (.A0(\rbzero.pov.ss_buffer[1] ),
    .A1(\rbzero.pov.ss_buffer[0] ),
    .S(_03084_),
    .X(_03552_));
 sky130_fd_sc_hd__clkbuf_1 _19880_ (.A(_03552_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _19881_ (.A0(net55),
    .A1(\rbzero.pov.sclk_buffer[0] ),
    .S(_09734_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_1 _19882_ (.A(_03553_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _19883_ (.A0(\rbzero.pov.sclk_buffer[1] ),
    .A1(\rbzero.pov.sclk_buffer[0] ),
    .S(_03084_),
    .X(_03554_));
 sky130_fd_sc_hd__clkbuf_1 _19884_ (.A(_03554_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _19885_ (.A0(\rbzero.pov.sclk_buffer[2] ),
    .A1(\rbzero.pov.sclk_buffer[1] ),
    .S(_08116_),
    .X(_03555_));
 sky130_fd_sc_hd__clkbuf_1 _19886_ (.A(_03555_),
    .X(_01166_));
 sky130_fd_sc_hd__nor2_1 _19887_ (.A(net41),
    .B(net40),
    .Y(_03556_));
 sky130_fd_sc_hd__and2_4 _19888_ (.A(\rbzero.pov.ready ),
    .B(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__o21ai_4 _19889_ (.A1(net40),
    .A2(_03557_),
    .B1(_03095_),
    .Y(_03558_));
 sky130_fd_sc_hd__clkbuf_4 _19890_ (.A(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__inv_2 _19891_ (.A(\rbzero.debug_overlay.playerX[-9] ),
    .Y(_03560_));
 sky130_fd_sc_hd__buf_4 _19892_ (.A(_03437_),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_1 _19893_ (.A0(_03560_),
    .A1(\rbzero.pov.ready_buffer[59] ),
    .S(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__nand2_1 _19894_ (.A(_03560_),
    .B(_03559_),
    .Y(_03563_));
 sky130_fd_sc_hd__o211a_1 _19895_ (.A1(_03559_),
    .A2(_03562_),
    .B1(_03563_),
    .C1(_03302_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _19896_ (.A0(_08186_),
    .A1(\rbzero.pov.ready_buffer[60] ),
    .S(_03561_),
    .X(_03564_));
 sky130_fd_sc_hd__o21a_2 _19897_ (.A1(net40),
    .A2(_03557_),
    .B1(_03095_),
    .X(_03565_));
 sky130_fd_sc_hd__or2_1 _19898_ (.A(\rbzero.debug_overlay.playerX[-8] ),
    .B(_03565_),
    .X(_03566_));
 sky130_fd_sc_hd__o211a_1 _19899_ (.A1(_03559_),
    .A2(_03564_),
    .B1(_03566_),
    .C1(_03302_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _19900_ (.A0(_08209_),
    .A1(\rbzero.pov.ready_buffer[61] ),
    .S(_03561_),
    .X(_03567_));
 sky130_fd_sc_hd__or2_1 _19901_ (.A(\rbzero.debug_overlay.playerX[-7] ),
    .B(_03565_),
    .X(_03568_));
 sky130_fd_sc_hd__o211a_1 _19902_ (.A1(_03559_),
    .A2(_03567_),
    .B1(_03568_),
    .C1(_03302_),
    .X(_01169_));
 sky130_fd_sc_hd__clkbuf_4 _19903_ (.A(_03565_),
    .X(_03569_));
 sky130_fd_sc_hd__buf_2 _19904_ (.A(_03437_),
    .X(_03570_));
 sky130_fd_sc_hd__nor2_1 _19905_ (.A(_08217_),
    .B(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__a211o_1 _19906_ (.A1(\rbzero.pov.ready_buffer[62] ),
    .A2(_03438_),
    .B1(_03559_),
    .C1(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__o211a_1 _19907_ (.A1(\rbzero.debug_overlay.playerX[-6] ),
    .A2(_03569_),
    .B1(_03572_),
    .C1(_03302_),
    .X(_01170_));
 sky130_fd_sc_hd__nor2_1 _19908_ (.A(_08239_),
    .B(_03570_),
    .Y(_03573_));
 sky130_fd_sc_hd__a211o_1 _19909_ (.A1(\rbzero.pov.ready_buffer[63] ),
    .A2(_03438_),
    .B1(_03558_),
    .C1(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__o211a_1 _19910_ (.A1(\rbzero.debug_overlay.playerX[-5] ),
    .A2(_03569_),
    .B1(_03574_),
    .C1(_03302_),
    .X(_01171_));
 sky130_fd_sc_hd__nor2_1 _19911_ (.A(_08256_),
    .B(_03570_),
    .Y(_03575_));
 sky130_fd_sc_hd__a211o_1 _19912_ (.A1(\rbzero.pov.ready_buffer[64] ),
    .A2(_03438_),
    .B1(_03558_),
    .C1(_03575_),
    .X(_03576_));
 sky130_fd_sc_hd__o211a_1 _19913_ (.A1(\rbzero.debug_overlay.playerX[-4] ),
    .A2(_03569_),
    .B1(_03576_),
    .C1(_03302_),
    .X(_01172_));
 sky130_fd_sc_hd__nor2_1 _19914_ (.A(_08279_),
    .B(_03570_),
    .Y(_03577_));
 sky130_fd_sc_hd__a211o_1 _19915_ (.A1(\rbzero.pov.ready_buffer[65] ),
    .A2(_03438_),
    .B1(_03558_),
    .C1(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__clkbuf_4 _19916_ (.A(_03212_),
    .X(_03579_));
 sky130_fd_sc_hd__o211a_1 _19917_ (.A1(\rbzero.debug_overlay.playerX[-3] ),
    .A2(_03569_),
    .B1(_03578_),
    .C1(_03579_),
    .X(_01173_));
 sky130_fd_sc_hd__nor2_1 _19918_ (.A(_08307_),
    .B(_03570_),
    .Y(_03580_));
 sky130_fd_sc_hd__a211o_1 _19919_ (.A1(\rbzero.pov.ready_buffer[66] ),
    .A2(_03438_),
    .B1(_03558_),
    .C1(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__o211a_1 _19920_ (.A1(\rbzero.debug_overlay.playerX[-2] ),
    .A2(_03569_),
    .B1(_03581_),
    .C1(_03579_),
    .X(_01174_));
 sky130_fd_sc_hd__nand2_1 _19921_ (.A(_03095_),
    .B(_03436_),
    .Y(_03582_));
 sky130_fd_sc_hd__o221a_1 _19922_ (.A1(\rbzero.pov.ready_buffer[67] ),
    .A2(_03436_),
    .B1(_03582_),
    .B2(_08317_),
    .C1(_03569_),
    .X(_03583_));
 sky130_fd_sc_hd__clkbuf_4 _19923_ (.A(_04409_),
    .X(_03584_));
 sky130_fd_sc_hd__a211o_1 _19924_ (.A1(\rbzero.debug_overlay.playerX[-1] ),
    .A2(_03559_),
    .B1(_03583_),
    .C1(_03584_),
    .X(_01175_));
 sky130_fd_sc_hd__nor2_1 _19925_ (.A(_03116_),
    .B(_03556_),
    .Y(_03585_));
 sky130_fd_sc_hd__buf_2 _19926_ (.A(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__or2_1 _19927_ (.A(\rbzero.debug_overlay.playerX[0] ),
    .B(_08315_),
    .X(_03587_));
 sky130_fd_sc_hd__inv_2 _19928_ (.A(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__a21o_1 _19929_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_08315_),
    .B1(_03582_),
    .X(_03589_));
 sky130_fd_sc_hd__o221a_1 _19930_ (.A1(\rbzero.pov.ready_buffer[68] ),
    .A2(_03586_),
    .B1(_03588_),
    .B2(_03589_),
    .C1(_03569_),
    .X(_03590_));
 sky130_fd_sc_hd__a211o_1 _19931_ (.A1(\rbzero.debug_overlay.playerX[0] ),
    .A2(_03559_),
    .B1(_03590_),
    .C1(_03584_),
    .X(_01176_));
 sky130_fd_sc_hd__nor2_1 _19932_ (.A(\rbzero.debug_overlay.playerX[1] ),
    .B(_03587_),
    .Y(_03591_));
 sky130_fd_sc_hd__a21o_1 _19933_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03587_),
    .B1(_03582_),
    .X(_03592_));
 sky130_fd_sc_hd__o221a_1 _19934_ (.A1(\rbzero.pov.ready_buffer[69] ),
    .A2(_03586_),
    .B1(_03591_),
    .B2(_03592_),
    .C1(_03569_),
    .X(_03593_));
 sky130_fd_sc_hd__a211o_1 _19935_ (.A1(\rbzero.debug_overlay.playerX[1] ),
    .A2(_03559_),
    .B1(_03593_),
    .C1(_03584_),
    .X(_01177_));
 sky130_fd_sc_hd__nand2_1 _19936_ (.A(_04674_),
    .B(_03591_),
    .Y(_03594_));
 sky130_fd_sc_hd__or2_1 _19937_ (.A(_04674_),
    .B(_03591_),
    .X(_03595_));
 sky130_fd_sc_hd__a21oi_1 _19938_ (.A1(_03594_),
    .A2(_03595_),
    .B1(_03561_),
    .Y(_03596_));
 sky130_fd_sc_hd__a211o_1 _19939_ (.A1(\rbzero.pov.ready_buffer[70] ),
    .A2(_03438_),
    .B1(_03558_),
    .C1(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__o211a_1 _19940_ (.A1(\rbzero.debug_overlay.playerX[2] ),
    .A2(_03569_),
    .B1(_03597_),
    .C1(_03579_),
    .X(_01178_));
 sky130_fd_sc_hd__or2_1 _19941_ (.A(\rbzero.debug_overlay.playerX[3] ),
    .B(_03594_),
    .X(_03598_));
 sky130_fd_sc_hd__and2_1 _19942_ (.A(_03436_),
    .B(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__inv_2 _19943_ (.A(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__a21o_1 _19944_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_03594_),
    .B1(_03116_),
    .X(_03601_));
 sky130_fd_sc_hd__o221a_1 _19945_ (.A1(\rbzero.pov.ready_buffer[71] ),
    .A2(_03586_),
    .B1(_03600_),
    .B2(_03601_),
    .C1(_03565_),
    .X(_03602_));
 sky130_fd_sc_hd__a211o_1 _19946_ (.A1(\rbzero.debug_overlay.playerX[3] ),
    .A2(_03559_),
    .B1(_03602_),
    .C1(_03584_),
    .X(_01179_));
 sky130_fd_sc_hd__o21a_1 _19947_ (.A1(_03559_),
    .A2(_03599_),
    .B1(\rbzero.debug_overlay.playerX[4] ),
    .X(_03603_));
 sky130_fd_sc_hd__nor2_1 _19948_ (.A(\rbzero.debug_overlay.playerX[4] ),
    .B(_03598_),
    .Y(_03604_));
 sky130_fd_sc_hd__o21a_1 _19949_ (.A1(_03556_),
    .A2(_03604_),
    .B1(_03565_),
    .X(_03605_));
 sky130_fd_sc_hd__o21a_1 _19950_ (.A1(\rbzero.pov.ready_buffer[72] ),
    .A2(_03586_),
    .B1(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__o21a_1 _19951_ (.A1(_03603_),
    .A2(_03606_),
    .B1(_03103_),
    .X(_01180_));
 sky130_fd_sc_hd__nor2_1 _19952_ (.A(_06133_),
    .B(_03605_),
    .Y(_03607_));
 sky130_fd_sc_hd__a21o_1 _19953_ (.A1(_06133_),
    .A2(_03604_),
    .B1(_03437_),
    .X(_03608_));
 sky130_fd_sc_hd__o211a_1 _19954_ (.A1(\rbzero.pov.ready_buffer[73] ),
    .A2(_03586_),
    .B1(_03569_),
    .C1(_03608_),
    .X(_03609_));
 sky130_fd_sc_hd__o21a_1 _19955_ (.A1(_03607_),
    .A2(_03609_),
    .B1(_03103_),
    .X(_01181_));
 sky130_fd_sc_hd__o21ai_4 _19956_ (.A1(net41),
    .A2(_03557_),
    .B1(_03095_),
    .Y(_03610_));
 sky130_fd_sc_hd__clkbuf_4 _19957_ (.A(_03610_),
    .X(_03611_));
 sky130_fd_sc_hd__mux2_1 _19958_ (.A0(_08437_),
    .A1(\rbzero.pov.ready_buffer[44] ),
    .S(_03561_),
    .X(_03612_));
 sky130_fd_sc_hd__nand2_1 _19959_ (.A(_08437_),
    .B(_03611_),
    .Y(_03613_));
 sky130_fd_sc_hd__o211a_1 _19960_ (.A1(_03611_),
    .A2(_03612_),
    .B1(_03613_),
    .C1(_03579_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _19961_ (.A0(_08189_),
    .A1(\rbzero.pov.ready_buffer[45] ),
    .S(_03561_),
    .X(_03614_));
 sky130_fd_sc_hd__nand2_1 _19962_ (.A(_08190_),
    .B(_03611_),
    .Y(_03615_));
 sky130_fd_sc_hd__o211a_1 _19963_ (.A1(_03611_),
    .A2(_03614_),
    .B1(_03615_),
    .C1(_03579_),
    .X(_01183_));
 sky130_fd_sc_hd__o21a_1 _19964_ (.A1(net41),
    .A2(_03557_),
    .B1(_03095_),
    .X(_03616_));
 sky130_fd_sc_hd__clkbuf_4 _19965_ (.A(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__nor2_1 _19966_ (.A(_08204_),
    .B(_03570_),
    .Y(_03618_));
 sky130_fd_sc_hd__a211o_1 _19967_ (.A1(\rbzero.pov.ready_buffer[46] ),
    .A2(_03438_),
    .B1(_03610_),
    .C1(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__o211a_1 _19968_ (.A1(\rbzero.debug_overlay.playerY[-7] ),
    .A2(_03617_),
    .B1(_03619_),
    .C1(_03579_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _19969_ (.A0(_08223_),
    .A1(\rbzero.pov.ready_buffer[47] ),
    .S(_03561_),
    .X(_03620_));
 sky130_fd_sc_hd__nand2_1 _19970_ (.A(_08220_),
    .B(_03611_),
    .Y(_03621_));
 sky130_fd_sc_hd__o211a_1 _19971_ (.A1(_03611_),
    .A2(_03620_),
    .B1(_03621_),
    .C1(_03579_),
    .X(_01185_));
 sky130_fd_sc_hd__nor2_1 _19972_ (.A(_08241_),
    .B(_03570_),
    .Y(_03622_));
 sky130_fd_sc_hd__a211o_1 _19973_ (.A1(\rbzero.pov.ready_buffer[48] ),
    .A2(_03438_),
    .B1(_03610_),
    .C1(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__o211a_1 _19974_ (.A1(\rbzero.debug_overlay.playerY[-5] ),
    .A2(_03617_),
    .B1(_03623_),
    .C1(_03579_),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _19975_ (.A0(_08261_),
    .A1(\rbzero.pov.ready_buffer[49] ),
    .S(_03561_),
    .X(_03624_));
 sky130_fd_sc_hd__nand2_1 _19976_ (.A(_08258_),
    .B(_03610_),
    .Y(_03625_));
 sky130_fd_sc_hd__o211a_1 _19977_ (.A1(_03611_),
    .A2(_03624_),
    .B1(_03625_),
    .C1(_03579_),
    .X(_01187_));
 sky130_fd_sc_hd__nor2_1 _19978_ (.A(_08283_),
    .B(_03570_),
    .Y(_03626_));
 sky130_fd_sc_hd__a211o_1 _19979_ (.A1(\rbzero.pov.ready_buffer[50] ),
    .A2(_03438_),
    .B1(_03610_),
    .C1(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__o211a_1 _19980_ (.A1(\rbzero.debug_overlay.playerY[-3] ),
    .A2(_03617_),
    .B1(_03627_),
    .C1(_03579_),
    .X(_01188_));
 sky130_fd_sc_hd__nor2_1 _19981_ (.A(_08309_),
    .B(_03561_),
    .Y(_03628_));
 sky130_fd_sc_hd__a211o_1 _19982_ (.A1(\rbzero.pov.ready_buffer[51] ),
    .A2(_03570_),
    .B1(_03610_),
    .C1(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__buf_4 _19983_ (.A(_03212_),
    .X(_03630_));
 sky130_fd_sc_hd__o211a_1 _19984_ (.A1(\rbzero.debug_overlay.playerY[-2] ),
    .A2(_03617_),
    .B1(_03629_),
    .C1(_03630_),
    .X(_01189_));
 sky130_fd_sc_hd__o221a_1 _19985_ (.A1(\rbzero.pov.ready_buffer[52] ),
    .A2(_03436_),
    .B1(_03582_),
    .B2(_08322_),
    .C1(_03617_),
    .X(_03631_));
 sky130_fd_sc_hd__a211o_1 _19986_ (.A1(\rbzero.debug_overlay.playerY[-1] ),
    .A2(_03611_),
    .B1(_03631_),
    .C1(_03584_),
    .X(_01190_));
 sky130_fd_sc_hd__or2_1 _19987_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_08320_),
    .X(_03632_));
 sky130_fd_sc_hd__nand2_1 _19988_ (.A(\rbzero.debug_overlay.playerY[0] ),
    .B(_08320_),
    .Y(_03633_));
 sky130_fd_sc_hd__a21oi_1 _19989_ (.A1(_03632_),
    .A2(_03633_),
    .B1(_03561_),
    .Y(_03634_));
 sky130_fd_sc_hd__a211o_1 _19990_ (.A1(\rbzero.pov.ready_buffer[53] ),
    .A2(_03570_),
    .B1(_03610_),
    .C1(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__o211a_1 _19991_ (.A1(\rbzero.debug_overlay.playerY[0] ),
    .A2(_03617_),
    .B1(_03635_),
    .C1(_03630_),
    .X(_01191_));
 sky130_fd_sc_hd__and2_1 _19992_ (.A(\rbzero.debug_overlay.playerY[1] ),
    .B(_03632_),
    .X(_03636_));
 sky130_fd_sc_hd__o21ai_1 _19993_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03632_),
    .B1(_03585_),
    .Y(_03637_));
 sky130_fd_sc_hd__o221a_1 _19994_ (.A1(\rbzero.pov.ready_buffer[54] ),
    .A2(_03586_),
    .B1(_03636_),
    .B2(_03637_),
    .C1(_03617_),
    .X(_03638_));
 sky130_fd_sc_hd__a211o_1 _19995_ (.A1(\rbzero.debug_overlay.playerY[1] ),
    .A2(_03611_),
    .B1(_03638_),
    .C1(_03584_),
    .X(_01192_));
 sky130_fd_sc_hd__a21o_1 _19996_ (.A1(_03617_),
    .A2(_03637_),
    .B1(_06112_),
    .X(_03639_));
 sky130_fd_sc_hd__or3_1 _19997_ (.A(\rbzero.debug_overlay.playerY[2] ),
    .B(\rbzero.debug_overlay.playerY[1] ),
    .C(_03632_),
    .X(_03640_));
 sky130_fd_sc_hd__nor2_1 _19998_ (.A(\rbzero.pov.ready_buffer[55] ),
    .B(_03585_),
    .Y(_03641_));
 sky130_fd_sc_hd__a211o_1 _19999_ (.A1(_03586_),
    .A2(_03640_),
    .B1(_03641_),
    .C1(_03610_),
    .X(_03642_));
 sky130_fd_sc_hd__a21oi_1 _20000_ (.A1(_03639_),
    .A2(_03642_),
    .B1(_03584_),
    .Y(_01193_));
 sky130_fd_sc_hd__o21a_1 _20001_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03640_),
    .B1(_03436_),
    .X(_03643_));
 sky130_fd_sc_hd__inv_2 _20002_ (.A(_03643_),
    .Y(_03644_));
 sky130_fd_sc_hd__a21o_1 _20003_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03640_),
    .B1(_03116_),
    .X(_03645_));
 sky130_fd_sc_hd__o221a_1 _20004_ (.A1(\rbzero.pov.ready_buffer[56] ),
    .A2(_03586_),
    .B1(_03644_),
    .B2(_03645_),
    .C1(_03617_),
    .X(_03646_));
 sky130_fd_sc_hd__a211o_1 _20005_ (.A1(\rbzero.debug_overlay.playerY[3] ),
    .A2(_03611_),
    .B1(_03646_),
    .C1(_03584_),
    .X(_01194_));
 sky130_fd_sc_hd__o21a_1 _20006_ (.A1(_03610_),
    .A2(_03643_),
    .B1(\rbzero.debug_overlay.playerY[4] ),
    .X(_03647_));
 sky130_fd_sc_hd__and3b_1 _20007_ (.A_N(_03640_),
    .B(_04667_),
    .C(_04673_),
    .X(_03648_));
 sky130_fd_sc_hd__o21a_1 _20008_ (.A1(_03556_),
    .A2(_03648_),
    .B1(_03616_),
    .X(_03649_));
 sky130_fd_sc_hd__o21a_1 _20009_ (.A1(\rbzero.pov.ready_buffer[57] ),
    .A2(_03586_),
    .B1(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__o21a_1 _20010_ (.A1(_03647_),
    .A2(_03650_),
    .B1(_03103_),
    .X(_01195_));
 sky130_fd_sc_hd__nor2_1 _20011_ (.A(_06114_),
    .B(_03649_),
    .Y(_03651_));
 sky130_fd_sc_hd__a21o_1 _20012_ (.A1(_06114_),
    .A2(_03648_),
    .B1(_03437_),
    .X(_03652_));
 sky130_fd_sc_hd__o211a_1 _20013_ (.A1(\rbzero.pov.ready_buffer[58] ),
    .A2(_03586_),
    .B1(_03617_),
    .C1(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__o21a_1 _20014_ (.A1(_03651_),
    .A2(_03653_),
    .B1(_03103_),
    .X(_01196_));
 sky130_fd_sc_hd__nand2_1 _20015_ (.A(_03095_),
    .B(_03557_),
    .Y(_03654_));
 sky130_fd_sc_hd__buf_2 _20016_ (.A(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__clkbuf_4 _20017_ (.A(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__and2_1 _20018_ (.A(_03095_),
    .B(_03557_),
    .X(_03657_));
 sky130_fd_sc_hd__buf_2 _20019_ (.A(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__or2_1 _20020_ (.A(\rbzero.debug_overlay.facingX[-9] ),
    .B(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__o211a_1 _20021_ (.A1(\rbzero.pov.ready_buffer[33] ),
    .A2(_03656_),
    .B1(_03659_),
    .C1(_03630_),
    .X(_01197_));
 sky130_fd_sc_hd__or2_1 _20022_ (.A(\rbzero.debug_overlay.facingX[-8] ),
    .B(_03658_),
    .X(_03660_));
 sky130_fd_sc_hd__o211a_1 _20023_ (.A1(\rbzero.pov.ready_buffer[34] ),
    .A2(_03656_),
    .B1(_03660_),
    .C1(_03630_),
    .X(_01198_));
 sky130_fd_sc_hd__or2_1 _20024_ (.A(\rbzero.debug_overlay.facingX[-7] ),
    .B(_03658_),
    .X(_03661_));
 sky130_fd_sc_hd__o211a_1 _20025_ (.A1(\rbzero.pov.ready_buffer[35] ),
    .A2(_03656_),
    .B1(_03661_),
    .C1(_03630_),
    .X(_01199_));
 sky130_fd_sc_hd__or2_1 _20026_ (.A(\rbzero.debug_overlay.facingX[-6] ),
    .B(_03658_),
    .X(_03662_));
 sky130_fd_sc_hd__o211a_1 _20027_ (.A1(\rbzero.pov.ready_buffer[36] ),
    .A2(_03656_),
    .B1(_03662_),
    .C1(_03630_),
    .X(_01200_));
 sky130_fd_sc_hd__clkbuf_4 _20028_ (.A(_03654_),
    .X(_03663_));
 sky130_fd_sc_hd__buf_2 _20029_ (.A(_03557_),
    .X(_03664_));
 sky130_fd_sc_hd__clkbuf_2 _20030_ (.A(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__and3_1 _20031_ (.A(\rbzero.pov.ready_buffer[37] ),
    .B(_03288_),
    .C(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__a211o_1 _20032_ (.A1(\rbzero.debug_overlay.facingX[-5] ),
    .A2(_03663_),
    .B1(_03666_),
    .C1(_03584_),
    .X(_01201_));
 sky130_fd_sc_hd__and3_1 _20033_ (.A(\rbzero.pov.ready_buffer[38] ),
    .B(_03288_),
    .C(_03665_),
    .X(_03667_));
 sky130_fd_sc_hd__a211o_1 _20034_ (.A1(\rbzero.debug_overlay.facingX[-4] ),
    .A2(_03663_),
    .B1(_03667_),
    .C1(_03584_),
    .X(_01202_));
 sky130_fd_sc_hd__and3_1 _20035_ (.A(\rbzero.pov.ready_buffer[39] ),
    .B(_03288_),
    .C(_03665_),
    .X(_03668_));
 sky130_fd_sc_hd__clkbuf_4 _20036_ (.A(_04409_),
    .X(_03669_));
 sky130_fd_sc_hd__a211o_1 _20037_ (.A1(\rbzero.debug_overlay.facingX[-3] ),
    .A2(_03663_),
    .B1(_03668_),
    .C1(_03669_),
    .X(_01203_));
 sky130_fd_sc_hd__or2_1 _20038_ (.A(\rbzero.debug_overlay.facingX[-2] ),
    .B(_03658_),
    .X(_03670_));
 sky130_fd_sc_hd__o211a_1 _20039_ (.A1(\rbzero.pov.ready_buffer[40] ),
    .A2(_03656_),
    .B1(_03670_),
    .C1(_03630_),
    .X(_01204_));
 sky130_fd_sc_hd__and3_1 _20040_ (.A(\rbzero.pov.ready_buffer[41] ),
    .B(_03288_),
    .C(_03665_),
    .X(_03671_));
 sky130_fd_sc_hd__a211o_1 _20041_ (.A1(\rbzero.debug_overlay.facingX[-1] ),
    .A2(_03663_),
    .B1(_03671_),
    .C1(_03669_),
    .X(_01205_));
 sky130_fd_sc_hd__or2_1 _20042_ (.A(\rbzero.debug_overlay.facingX[0] ),
    .B(_03658_),
    .X(_03672_));
 sky130_fd_sc_hd__o211a_1 _20043_ (.A1(\rbzero.pov.ready_buffer[42] ),
    .A2(_03656_),
    .B1(_03672_),
    .C1(_03630_),
    .X(_01206_));
 sky130_fd_sc_hd__or2_1 _20044_ (.A(\rbzero.debug_overlay.facingX[10] ),
    .B(_03658_),
    .X(_03673_));
 sky130_fd_sc_hd__o211a_1 _20045_ (.A1(net512),
    .A2(_03656_),
    .B1(_03673_),
    .C1(_03630_),
    .X(_01207_));
 sky130_fd_sc_hd__and3_1 _20046_ (.A(\rbzero.pov.ready_buffer[22] ),
    .B(_03288_),
    .C(_03665_),
    .X(_03674_));
 sky130_fd_sc_hd__a211o_1 _20047_ (.A1(\rbzero.debug_overlay.facingY[-9] ),
    .A2(_03663_),
    .B1(_03674_),
    .C1(_03669_),
    .X(_01208_));
 sky130_fd_sc_hd__or2_1 _20048_ (.A(\rbzero.debug_overlay.facingY[-8] ),
    .B(_03658_),
    .X(_03675_));
 sky130_fd_sc_hd__o211a_1 _20049_ (.A1(\rbzero.pov.ready_buffer[23] ),
    .A2(_03656_),
    .B1(_03675_),
    .C1(_03630_),
    .X(_01209_));
 sky130_fd_sc_hd__clkbuf_4 _20050_ (.A(_03654_),
    .X(_03676_));
 sky130_fd_sc_hd__and3_1 _20051_ (.A(\rbzero.pov.ready_buffer[24] ),
    .B(_03288_),
    .C(_03665_),
    .X(_03677_));
 sky130_fd_sc_hd__a211o_1 _20052_ (.A1(\rbzero.debug_overlay.facingY[-7] ),
    .A2(_03676_),
    .B1(_03677_),
    .C1(_03669_),
    .X(_01210_));
 sky130_fd_sc_hd__and3_1 _20053_ (.A(\rbzero.pov.ready_buffer[25] ),
    .B(_03288_),
    .C(_03665_),
    .X(_03678_));
 sky130_fd_sc_hd__a211o_1 _20054_ (.A1(\rbzero.debug_overlay.facingY[-6] ),
    .A2(_03676_),
    .B1(_03678_),
    .C1(_03669_),
    .X(_01211_));
 sky130_fd_sc_hd__and3_1 _20055_ (.A(\rbzero.pov.ready_buffer[26] ),
    .B(_03288_),
    .C(_03665_),
    .X(_03679_));
 sky130_fd_sc_hd__a211o_1 _20056_ (.A1(\rbzero.debug_overlay.facingY[-5] ),
    .A2(_03676_),
    .B1(_03679_),
    .C1(_03669_),
    .X(_01212_));
 sky130_fd_sc_hd__or2_1 _20057_ (.A(\rbzero.debug_overlay.facingY[-4] ),
    .B(_03658_),
    .X(_03680_));
 sky130_fd_sc_hd__clkbuf_4 _20058_ (.A(_03212_),
    .X(_03681_));
 sky130_fd_sc_hd__o211a_1 _20059_ (.A1(\rbzero.pov.ready_buffer[27] ),
    .A2(_03656_),
    .B1(_03680_),
    .C1(_03681_),
    .X(_01213_));
 sky130_fd_sc_hd__or2_1 _20060_ (.A(\rbzero.debug_overlay.facingY[-3] ),
    .B(_03658_),
    .X(_03682_));
 sky130_fd_sc_hd__o211a_1 _20061_ (.A1(\rbzero.pov.ready_buffer[28] ),
    .A2(_03656_),
    .B1(_03682_),
    .C1(_03681_),
    .X(_01214_));
 sky130_fd_sc_hd__and3_1 _20062_ (.A(\rbzero.pov.ready_buffer[29] ),
    .B(_03288_),
    .C(_03665_),
    .X(_03683_));
 sky130_fd_sc_hd__a211o_1 _20063_ (.A1(\rbzero.debug_overlay.facingY[-2] ),
    .A2(_03676_),
    .B1(_03683_),
    .C1(_03669_),
    .X(_01215_));
 sky130_fd_sc_hd__clkbuf_4 _20064_ (.A(_03654_),
    .X(_03684_));
 sky130_fd_sc_hd__buf_2 _20065_ (.A(_03657_),
    .X(_03685_));
 sky130_fd_sc_hd__or2_1 _20066_ (.A(\rbzero.debug_overlay.facingY[-1] ),
    .B(_03685_),
    .X(_03686_));
 sky130_fd_sc_hd__o211a_1 _20067_ (.A1(\rbzero.pov.ready_buffer[30] ),
    .A2(_03684_),
    .B1(_03686_),
    .C1(_03681_),
    .X(_01216_));
 sky130_fd_sc_hd__buf_2 _20068_ (.A(_03096_),
    .X(_03687_));
 sky130_fd_sc_hd__and3_1 _20069_ (.A(\rbzero.pov.ready_buffer[31] ),
    .B(_03687_),
    .C(_03665_),
    .X(_03688_));
 sky130_fd_sc_hd__a211o_1 _20070_ (.A1(\rbzero.debug_overlay.facingY[0] ),
    .A2(_03676_),
    .B1(_03688_),
    .C1(_03669_),
    .X(_01217_));
 sky130_fd_sc_hd__and3_1 _20071_ (.A(\rbzero.pov.ready_buffer[32] ),
    .B(_03687_),
    .C(_03664_),
    .X(_03689_));
 sky130_fd_sc_hd__a211o_1 _20072_ (.A1(\rbzero.debug_overlay.facingY[10] ),
    .A2(_03676_),
    .B1(_03689_),
    .C1(_03669_),
    .X(_01218_));
 sky130_fd_sc_hd__and3_1 _20073_ (.A(\rbzero.pov.ready_buffer[11] ),
    .B(_03687_),
    .C(_03664_),
    .X(_03690_));
 sky130_fd_sc_hd__a211o_1 _20074_ (.A1(\rbzero.debug_overlay.vplaneX[-9] ),
    .A2(_03676_),
    .B1(_03690_),
    .C1(_03669_),
    .X(_01219_));
 sky130_fd_sc_hd__or2_1 _20075_ (.A(\rbzero.debug_overlay.vplaneX[-8] ),
    .B(_03685_),
    .X(_03691_));
 sky130_fd_sc_hd__o211a_1 _20076_ (.A1(\rbzero.pov.ready_buffer[12] ),
    .A2(_03684_),
    .B1(_03691_),
    .C1(_03681_),
    .X(_01220_));
 sky130_fd_sc_hd__or2_1 _20077_ (.A(\rbzero.debug_overlay.vplaneX[-7] ),
    .B(_03685_),
    .X(_03692_));
 sky130_fd_sc_hd__o211a_1 _20078_ (.A1(\rbzero.pov.ready_buffer[13] ),
    .A2(_03684_),
    .B1(_03692_),
    .C1(_03681_),
    .X(_01221_));
 sky130_fd_sc_hd__or2_1 _20079_ (.A(_05120_),
    .B(_03685_),
    .X(_03693_));
 sky130_fd_sc_hd__o211a_1 _20080_ (.A1(\rbzero.pov.ready_buffer[14] ),
    .A2(_03684_),
    .B1(_03693_),
    .C1(_03681_),
    .X(_01222_));
 sky130_fd_sc_hd__and3_1 _20081_ (.A(\rbzero.pov.ready_buffer[15] ),
    .B(_03687_),
    .C(_03664_),
    .X(_03694_));
 sky130_fd_sc_hd__buf_4 _20082_ (.A(_09734_),
    .X(_03695_));
 sky130_fd_sc_hd__a211o_1 _20083_ (.A1(_05111_),
    .A2(_03676_),
    .B1(_03694_),
    .C1(_03695_),
    .X(_01223_));
 sky130_fd_sc_hd__and3_1 _20084_ (.A(\rbzero.pov.ready_buffer[16] ),
    .B(_03687_),
    .C(_03664_),
    .X(_03696_));
 sky130_fd_sc_hd__a211o_1 _20085_ (.A1(\rbzero.debug_overlay.vplaneX[-4] ),
    .A2(_03676_),
    .B1(_03696_),
    .C1(_03695_),
    .X(_01224_));
 sky130_fd_sc_hd__or2_1 _20086_ (.A(\rbzero.debug_overlay.vplaneX[-3] ),
    .B(_03685_),
    .X(_03697_));
 sky130_fd_sc_hd__o211a_1 _20087_ (.A1(\rbzero.pov.ready_buffer[17] ),
    .A2(_03684_),
    .B1(_03697_),
    .C1(_03681_),
    .X(_01225_));
 sky130_fd_sc_hd__and3_1 _20088_ (.A(\rbzero.pov.ready_buffer[18] ),
    .B(_03687_),
    .C(_03664_),
    .X(_03698_));
 sky130_fd_sc_hd__a211o_1 _20089_ (.A1(_05106_),
    .A2(_03676_),
    .B1(_03698_),
    .C1(_03695_),
    .X(_01226_));
 sky130_fd_sc_hd__or2_1 _20090_ (.A(\rbzero.debug_overlay.vplaneX[-1] ),
    .B(_03685_),
    .X(_03699_));
 sky130_fd_sc_hd__o211a_1 _20091_ (.A1(\rbzero.pov.ready_buffer[19] ),
    .A2(_03684_),
    .B1(_03699_),
    .C1(_03681_),
    .X(_01227_));
 sky130_fd_sc_hd__nand2_1 _20092_ (.A(_02681_),
    .B(_03655_),
    .Y(_03700_));
 sky130_fd_sc_hd__o211a_1 _20093_ (.A1(\rbzero.pov.ready_buffer[20] ),
    .A2(_03684_),
    .B1(_03700_),
    .C1(_03681_),
    .X(_01228_));
 sky130_fd_sc_hd__nand2_1 _20094_ (.A(_02694_),
    .B(_03655_),
    .Y(_03701_));
 sky130_fd_sc_hd__o211a_1 _20095_ (.A1(\rbzero.pov.ready_buffer[21] ),
    .A2(_03684_),
    .B1(_03701_),
    .C1(_03681_),
    .X(_01229_));
 sky130_fd_sc_hd__nand2_1 _20096_ (.A(_02756_),
    .B(_03655_),
    .Y(_03702_));
 sky130_fd_sc_hd__buf_4 _20097_ (.A(_03084_),
    .X(_03703_));
 sky130_fd_sc_hd__o211a_1 _20098_ (.A1(\rbzero.pov.ready_buffer[0] ),
    .A2(_03684_),
    .B1(_03702_),
    .C1(_03703_),
    .X(_01230_));
 sky130_fd_sc_hd__or2_1 _20099_ (.A(\rbzero.debug_overlay.vplaneY[-8] ),
    .B(_03685_),
    .X(_03704_));
 sky130_fd_sc_hd__o211a_1 _20100_ (.A1(\rbzero.pov.ready_buffer[1] ),
    .A2(_03684_),
    .B1(_03704_),
    .C1(_03703_),
    .X(_01231_));
 sky130_fd_sc_hd__or2_1 _20101_ (.A(\rbzero.debug_overlay.vplaneY[-7] ),
    .B(_03685_),
    .X(_03705_));
 sky130_fd_sc_hd__o211a_1 _20102_ (.A1(\rbzero.pov.ready_buffer[2] ),
    .A2(_03663_),
    .B1(_03705_),
    .C1(_03703_),
    .X(_01232_));
 sky130_fd_sc_hd__and3_1 _20103_ (.A(\rbzero.pov.ready_buffer[3] ),
    .B(_03687_),
    .C(_03664_),
    .X(_03706_));
 sky130_fd_sc_hd__a211o_1 _20104_ (.A1(_05129_),
    .A2(_03655_),
    .B1(_03706_),
    .C1(_03695_),
    .X(_01233_));
 sky130_fd_sc_hd__and3_1 _20105_ (.A(\rbzero.pov.ready_buffer[4] ),
    .B(_03687_),
    .C(_03664_),
    .X(_03707_));
 sky130_fd_sc_hd__a211o_1 _20106_ (.A1(\rbzero.debug_overlay.vplaneY[-5] ),
    .A2(_03655_),
    .B1(_03707_),
    .C1(_03695_),
    .X(_01234_));
 sky130_fd_sc_hd__and3_1 _20107_ (.A(\rbzero.pov.ready_buffer[5] ),
    .B(_03687_),
    .C(_03664_),
    .X(_03708_));
 sky130_fd_sc_hd__a211o_1 _20108_ (.A1(_05132_),
    .A2(_03655_),
    .B1(_03708_),
    .C1(_03695_),
    .X(_01235_));
 sky130_fd_sc_hd__or2_1 _20109_ (.A(\rbzero.debug_overlay.vplaneY[-3] ),
    .B(_03685_),
    .X(_03709_));
 sky130_fd_sc_hd__o211a_1 _20110_ (.A1(\rbzero.pov.ready_buffer[6] ),
    .A2(_03663_),
    .B1(_03709_),
    .C1(_03703_),
    .X(_01236_));
 sky130_fd_sc_hd__and3_1 _20111_ (.A(\rbzero.pov.ready_buffer[7] ),
    .B(_03687_),
    .C(_03664_),
    .X(_03710_));
 sky130_fd_sc_hd__a211o_1 _20112_ (.A1(\rbzero.debug_overlay.vplaneY[-2] ),
    .A2(_03655_),
    .B1(_03710_),
    .C1(_03695_),
    .X(_01237_));
 sky130_fd_sc_hd__or2_1 _20113_ (.A(\rbzero.debug_overlay.vplaneY[-1] ),
    .B(_03685_),
    .X(_03711_));
 sky130_fd_sc_hd__o211a_1 _20114_ (.A1(\rbzero.pov.ready_buffer[8] ),
    .A2(_03663_),
    .B1(_03711_),
    .C1(_03703_),
    .X(_01238_));
 sky130_fd_sc_hd__nand2_1 _20115_ (.A(_02907_),
    .B(_03655_),
    .Y(_03712_));
 sky130_fd_sc_hd__o211a_1 _20116_ (.A1(\rbzero.pov.ready_buffer[9] ),
    .A2(_03663_),
    .B1(_03712_),
    .C1(_03703_),
    .X(_01239_));
 sky130_fd_sc_hd__nand2_1 _20117_ (.A(_02889_),
    .B(_03655_),
    .Y(_03713_));
 sky130_fd_sc_hd__o211a_1 _20118_ (.A1(\rbzero.pov.ready_buffer[10] ),
    .A2(_03663_),
    .B1(_03713_),
    .C1(_03703_),
    .X(_01240_));
 sky130_fd_sc_hd__a31o_1 _20119_ (.A1(_03440_),
    .A2(_03439_),
    .A3(_03445_),
    .B1(\rbzero.pov.spi_done ),
    .X(_03714_));
 sky130_fd_sc_hd__and2_1 _20120_ (.A(_02968_),
    .B(_03714_),
    .X(_03715_));
 sky130_fd_sc_hd__clkbuf_1 _20121_ (.A(_03715_),
    .X(_01241_));
 sky130_fd_sc_hd__inv_2 _20122_ (.A(_04687_),
    .Y(_03716_));
 sky130_fd_sc_hd__and4b_1 _20123_ (.A_N(_05648_),
    .B(_05651_),
    .C(_03091_),
    .D(_04657_),
    .X(_03717_));
 sky130_fd_sc_hd__and4_1 _20124_ (.A(_05644_),
    .B(_03716_),
    .C(_04691_),
    .D(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__or4bb_1 _20125_ (.A(_05651_),
    .B(_05650_),
    .C_N(_05644_),
    .D_N(_04687_),
    .X(_03719_));
 sky130_fd_sc_hd__or4b_1 _20126_ (.A(_04731_),
    .B(_03719_),
    .C(_05648_),
    .D_N(_03091_),
    .X(_03720_));
 sky130_fd_sc_hd__o211a_1 _20127_ (.A1(\rbzero.vga_sync.vsync ),
    .A2(_03718_),
    .B1(_03720_),
    .C1(_03703_),
    .X(_01242_));
 sky130_fd_sc_hd__and3b_1 _20128_ (.A_N(_04698_),
    .B(_04413_),
    .C(_03977_),
    .X(_03721_));
 sky130_fd_sc_hd__a31o_1 _20129_ (.A1(_04589_),
    .A2(_05283_),
    .A3(_03721_),
    .B1(_04408_),
    .X(_03722_));
 sky130_fd_sc_hd__a31o_1 _20130_ (.A1(_03973_),
    .A2(_09727_),
    .A3(_03721_),
    .B1(\rbzero.hsync ),
    .X(_03723_));
 sky130_fd_sc_hd__and2b_1 _20131_ (.A_N(_03722_),
    .B(_03723_),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_1 _20132_ (.A(_03724_),
    .X(_01243_));
 sky130_fd_sc_hd__or4b_1 _20133_ (.A(_05652_),
    .B(_04695_),
    .C(_03719_),
    .D_N(_05653_),
    .X(_03725_));
 sky130_fd_sc_hd__and2_1 _20134_ (.A(_09729_),
    .B(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__nand2_1 _20135_ (.A(_05650_),
    .B(_09729_),
    .Y(_03727_));
 sky130_fd_sc_hd__o211a_1 _20136_ (.A1(_05650_),
    .A2(_03726_),
    .B1(_03727_),
    .C1(_03703_),
    .X(_01244_));
 sky130_fd_sc_hd__clkbuf_4 _20137_ (.A(_08116_),
    .X(_03728_));
 sky130_fd_sc_hd__nand3_1 _20138_ (.A(_05651_),
    .B(_05650_),
    .C(_09729_),
    .Y(_03729_));
 sky130_fd_sc_hd__a21o_1 _20139_ (.A1(_05650_),
    .A2(_09729_),
    .B1(_05651_),
    .X(_03730_));
 sky130_fd_sc_hd__and3_1 _20140_ (.A(_03728_),
    .B(_03729_),
    .C(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__clkbuf_1 _20141_ (.A(_03731_),
    .X(_01245_));
 sky130_fd_sc_hd__a21o_1 _20142_ (.A1(_08116_),
    .A2(_03725_),
    .B1(_09731_),
    .X(_03732_));
 sky130_fd_sc_hd__a21bo_1 _20143_ (.A1(_09729_),
    .A2(_03092_),
    .B1_N(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__a21oi_1 _20144_ (.A1(_03716_),
    .A2(_03729_),
    .B1(_03733_),
    .Y(_01246_));
 sky130_fd_sc_hd__buf_4 _20145_ (.A(_09732_),
    .X(_03734_));
 sky130_fd_sc_hd__a21oi_1 _20146_ (.A1(_05644_),
    .A2(_03092_),
    .B1(_04408_),
    .Y(_03735_));
 sky130_fd_sc_hd__o21a_1 _20147_ (.A1(_05644_),
    .A2(_03092_),
    .B1(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__a22o_1 _20148_ (.A1(_05644_),
    .A2(_03734_),
    .B1(_03726_),
    .B2(_03736_),
    .X(_01247_));
 sky130_fd_sc_hd__and2_1 _20149_ (.A(_05648_),
    .B(_03093_),
    .X(_03737_));
 sky130_fd_sc_hd__inv_2 _20150_ (.A(_03737_),
    .Y(_03738_));
 sky130_fd_sc_hd__o211a_1 _20151_ (.A1(_05648_),
    .A2(_03099_),
    .B1(_03738_),
    .C1(_03703_),
    .X(_01248_));
 sky130_fd_sc_hd__and3_1 _20152_ (.A(_04657_),
    .B(_05648_),
    .C(_03099_),
    .X(_03739_));
 sky130_fd_sc_hd__buf_4 _20153_ (.A(_09734_),
    .X(_03740_));
 sky130_fd_sc_hd__a211oi_1 _20154_ (.A1(_04731_),
    .A2(_03738_),
    .B1(_03739_),
    .C1(_03740_),
    .Y(_01249_));
 sky130_fd_sc_hd__nor2_1 _20155_ (.A(_04731_),
    .B(_03738_),
    .Y(_03741_));
 sky130_fd_sc_hd__nand2_1 _20156_ (.A(_05645_),
    .B(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__o211a_1 _20157_ (.A1(_05645_),
    .A2(_03739_),
    .B1(_03742_),
    .C1(_03118_),
    .X(_01250_));
 sky130_fd_sc_hd__nand2_1 _20158_ (.A(_04670_),
    .B(_03742_),
    .Y(_03743_));
 sky130_fd_sc_hd__nand2_1 _20159_ (.A(_05054_),
    .B(_03737_),
    .Y(_03744_));
 sky130_fd_sc_hd__and3_1 _20160_ (.A(_03728_),
    .B(_03743_),
    .C(_03744_),
    .X(_03745_));
 sky130_fd_sc_hd__clkbuf_1 _20161_ (.A(_03745_),
    .X(_01251_));
 sky130_fd_sc_hd__inv_2 _20162_ (.A(_05652_),
    .Y(_03746_));
 sky130_fd_sc_hd__and4_1 _20163_ (.A(_05652_),
    .B(_04642_),
    .C(_05645_),
    .D(_03741_),
    .X(_03747_));
 sky130_fd_sc_hd__a211oi_1 _20164_ (.A1(_03746_),
    .A2(_03744_),
    .B1(_03747_),
    .C1(_04409_),
    .Y(_01252_));
 sky130_fd_sc_hd__or2_1 _20165_ (.A(_05653_),
    .B(_03747_),
    .X(_03748_));
 sky130_fd_sc_hd__nand2_1 _20166_ (.A(_05653_),
    .B(_03747_),
    .Y(_03749_));
 sky130_fd_sc_hd__and3_1 _20167_ (.A(_03732_),
    .B(_03748_),
    .C(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__clkbuf_1 _20168_ (.A(_03750_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _20169_ (.A0(\rbzero.spi_registers.new_texadd[3][0] ),
    .A1(\rbzero.spi_registers.spi_buffer[0] ),
    .S(_03385_),
    .X(_03751_));
 sky130_fd_sc_hd__clkbuf_1 _20170_ (.A(_03751_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _20171_ (.A0(\rbzero.spi_registers.new_texadd[3][1] ),
    .A1(\rbzero.spi_registers.spi_buffer[1] ),
    .S(_03385_),
    .X(_03752_));
 sky130_fd_sc_hd__clkbuf_1 _20172_ (.A(_03752_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _20173_ (.A0(\rbzero.spi_registers.new_texadd[3][2] ),
    .A1(\rbzero.spi_registers.spi_buffer[2] ),
    .S(_03385_),
    .X(_03753_));
 sky130_fd_sc_hd__clkbuf_1 _20174_ (.A(_03753_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _20175_ (.A0(\rbzero.spi_registers.new_texadd[3][3] ),
    .A1(\rbzero.spi_registers.spi_buffer[3] ),
    .S(_03385_),
    .X(_03754_));
 sky130_fd_sc_hd__clkbuf_1 _20176_ (.A(_03754_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _20177_ (.A0(\rbzero.spi_registers.new_texadd[3][4] ),
    .A1(\rbzero.spi_registers.spi_buffer[4] ),
    .S(_03385_),
    .X(_03755_));
 sky130_fd_sc_hd__clkbuf_1 _20178_ (.A(_03755_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _20179_ (.A0(\rbzero.spi_registers.new_texadd[3][5] ),
    .A1(\rbzero.spi_registers.spi_buffer[5] ),
    .S(_03385_),
    .X(_03756_));
 sky130_fd_sc_hd__clkbuf_1 _20180_ (.A(_03756_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _20181_ (.A0(\rbzero.spi_registers.new_texadd[3][6] ),
    .A1(\rbzero.spi_registers.spi_buffer[6] ),
    .S(_03385_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_1 _20182_ (.A(_03757_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _20183_ (.A0(\rbzero.spi_registers.new_texadd[3][7] ),
    .A1(\rbzero.spi_registers.spi_buffer[7] ),
    .S(_03385_),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_1 _20184_ (.A(_03758_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _20185_ (.A0(\rbzero.spi_registers.new_texadd[3][8] ),
    .A1(\rbzero.spi_registers.spi_buffer[8] ),
    .S(_03385_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_1 _20186_ (.A(_03759_),
    .X(_01262_));
 sky130_fd_sc_hd__buf_4 _20187_ (.A(_03384_),
    .X(_03760_));
 sky130_fd_sc_hd__mux2_1 _20188_ (.A0(\rbzero.spi_registers.new_texadd[3][9] ),
    .A1(\rbzero.spi_registers.spi_buffer[9] ),
    .S(_03760_),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_1 _20189_ (.A(_03761_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _20190_ (.A0(\rbzero.spi_registers.new_texadd[3][10] ),
    .A1(\rbzero.spi_registers.spi_buffer[10] ),
    .S(_03760_),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_1 _20191_ (.A(_03762_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _20192_ (.A0(\rbzero.spi_registers.new_texadd[3][11] ),
    .A1(\rbzero.spi_registers.spi_buffer[11] ),
    .S(_03760_),
    .X(_03763_));
 sky130_fd_sc_hd__clkbuf_1 _20193_ (.A(_03763_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _20194_ (.A0(\rbzero.spi_registers.new_texadd[3][12] ),
    .A1(\rbzero.spi_registers.spi_buffer[12] ),
    .S(_03760_),
    .X(_03764_));
 sky130_fd_sc_hd__clkbuf_1 _20195_ (.A(_03764_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _20196_ (.A0(\rbzero.spi_registers.new_texadd[3][13] ),
    .A1(\rbzero.spi_registers.spi_buffer[13] ),
    .S(_03760_),
    .X(_03765_));
 sky130_fd_sc_hd__clkbuf_1 _20197_ (.A(_03765_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _20198_ (.A0(\rbzero.spi_registers.new_texadd[3][14] ),
    .A1(\rbzero.spi_registers.spi_buffer[14] ),
    .S(_03760_),
    .X(_03766_));
 sky130_fd_sc_hd__clkbuf_1 _20199_ (.A(_03766_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _20200_ (.A0(\rbzero.spi_registers.new_texadd[3][15] ),
    .A1(\rbzero.spi_registers.spi_buffer[15] ),
    .S(_03760_),
    .X(_03767_));
 sky130_fd_sc_hd__clkbuf_1 _20201_ (.A(_03767_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _20202_ (.A0(\rbzero.spi_registers.new_texadd[3][16] ),
    .A1(\rbzero.spi_registers.spi_buffer[16] ),
    .S(_03760_),
    .X(_03768_));
 sky130_fd_sc_hd__clkbuf_1 _20203_ (.A(_03768_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _20204_ (.A0(\rbzero.spi_registers.new_texadd[3][17] ),
    .A1(\rbzero.spi_registers.spi_buffer[17] ),
    .S(_03760_),
    .X(_03769_));
 sky130_fd_sc_hd__clkbuf_1 _20205_ (.A(_03769_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _20206_ (.A0(\rbzero.spi_registers.new_texadd[3][18] ),
    .A1(\rbzero.spi_registers.spi_buffer[18] ),
    .S(_03760_),
    .X(_03770_));
 sky130_fd_sc_hd__clkbuf_1 _20207_ (.A(_03770_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _20208_ (.A0(\rbzero.spi_registers.new_texadd[3][19] ),
    .A1(\rbzero.spi_registers.spi_buffer[19] ),
    .S(_03384_),
    .X(_03771_));
 sky130_fd_sc_hd__clkbuf_1 _20209_ (.A(_03771_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _20210_ (.A0(\rbzero.spi_registers.new_texadd[3][20] ),
    .A1(\rbzero.spi_registers.spi_buffer[20] ),
    .S(_03384_),
    .X(_03772_));
 sky130_fd_sc_hd__clkbuf_1 _20211_ (.A(_03772_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _20212_ (.A0(\rbzero.spi_registers.new_texadd[3][21] ),
    .A1(\rbzero.spi_registers.spi_buffer[21] ),
    .S(_03384_),
    .X(_03773_));
 sky130_fd_sc_hd__clkbuf_1 _20213_ (.A(_03773_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _20214_ (.A0(\rbzero.spi_registers.new_texadd[3][22] ),
    .A1(\rbzero.spi_registers.spi_buffer[22] ),
    .S(_03384_),
    .X(_03774_));
 sky130_fd_sc_hd__clkbuf_1 _20215_ (.A(_03774_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _20216_ (.A0(\rbzero.spi_registers.new_texadd[3][23] ),
    .A1(\rbzero.spi_registers.spi_buffer[23] ),
    .S(_03384_),
    .X(_03775_));
 sky130_fd_sc_hd__clkbuf_1 _20217_ (.A(_03775_),
    .X(_01277_));
 sky130_fd_sc_hd__inv_2 _20219__92 (.A(clknet_1_1__leaf__03465_),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _20220__93 (.A(clknet_1_1__leaf__03465_),
    .Y(net217));
 sky130_fd_sc_hd__inv_2 _20221__94 (.A(clknet_1_1__leaf__03465_),
    .Y(net218));
 sky130_fd_sc_hd__inv_2 _20222__95 (.A(clknet_1_1__leaf__03465_),
    .Y(net219));
 sky130_fd_sc_hd__inv_2 _20223__96 (.A(clknet_1_1__leaf__03465_),
    .Y(net220));
 sky130_fd_sc_hd__inv_2 _20225__97 (.A(clknet_1_0__leaf__03776_),
    .Y(net221));
 sky130_fd_sc_hd__buf_1 _20224_ (.A(clknet_1_0__leaf__03464_),
    .X(_03776_));
 sky130_fd_sc_hd__inv_2 _20226__98 (.A(clknet_1_0__leaf__03776_),
    .Y(net222));
 sky130_fd_sc_hd__inv_2 _20227__99 (.A(clknet_1_0__leaf__03776_),
    .Y(net223));
 sky130_fd_sc_hd__inv_2 _20228__100 (.A(clknet_1_0__leaf__03776_),
    .Y(net224));
 sky130_fd_sc_hd__inv_2 _20229__101 (.A(clknet_1_1__leaf__03776_),
    .Y(net225));
 sky130_fd_sc_hd__inv_2 _20230__102 (.A(clknet_1_1__leaf__03776_),
    .Y(net226));
 sky130_fd_sc_hd__inv_2 _20231__103 (.A(clknet_1_1__leaf__03776_),
    .Y(net227));
 sky130_fd_sc_hd__inv_2 _20232__104 (.A(clknet_1_1__leaf__03776_),
    .Y(net228));
 sky130_fd_sc_hd__inv_2 _20233__105 (.A(clknet_1_1__leaf__03776_),
    .Y(net229));
 sky130_fd_sc_hd__inv_2 _20234__106 (.A(clknet_1_1__leaf__03776_),
    .Y(net230));
 sky130_fd_sc_hd__inv_2 _20236__107 (.A(clknet_1_1__leaf__03777_),
    .Y(net231));
 sky130_fd_sc_hd__buf_1 _20235_ (.A(clknet_1_0__leaf__03464_),
    .X(_03777_));
 sky130_fd_sc_hd__inv_2 _20237__108 (.A(clknet_1_1__leaf__03777_),
    .Y(net232));
 sky130_fd_sc_hd__inv_2 _20238__109 (.A(clknet_1_0__leaf__03777_),
    .Y(net233));
 sky130_fd_sc_hd__inv_2 _20239__110 (.A(clknet_1_1__leaf__03777_),
    .Y(net234));
 sky130_fd_sc_hd__inv_2 _20240__111 (.A(clknet_1_1__leaf__03777_),
    .Y(net235));
 sky130_fd_sc_hd__inv_2 _20241__112 (.A(clknet_1_1__leaf__03777_),
    .Y(net236));
 sky130_fd_sc_hd__inv_2 _20242__113 (.A(clknet_1_1__leaf__03777_),
    .Y(net237));
 sky130_fd_sc_hd__inv_2 _20243__114 (.A(clknet_1_0__leaf__03777_),
    .Y(net238));
 sky130_fd_sc_hd__inv_2 _20244__115 (.A(clknet_1_0__leaf__03777_),
    .Y(net239));
 sky130_fd_sc_hd__inv_2 _20245__116 (.A(clknet_1_0__leaf__03777_),
    .Y(net240));
 sky130_fd_sc_hd__inv_2 _20247__117 (.A(clknet_1_0__leaf__03778_),
    .Y(net241));
 sky130_fd_sc_hd__buf_1 _20246_ (.A(clknet_1_0__leaf__03464_),
    .X(_03778_));
 sky130_fd_sc_hd__inv_2 _20248__118 (.A(clknet_1_0__leaf__03778_),
    .Y(net242));
 sky130_fd_sc_hd__inv_2 _20249__119 (.A(clknet_1_0__leaf__03778_),
    .Y(net243));
 sky130_fd_sc_hd__inv_2 _20250__120 (.A(clknet_1_0__leaf__03778_),
    .Y(net244));
 sky130_fd_sc_hd__inv_2 _20251__121 (.A(clknet_1_1__leaf__03778_),
    .Y(net245));
 sky130_fd_sc_hd__inv_2 _20252__122 (.A(clknet_1_0__leaf__03778_),
    .Y(net246));
 sky130_fd_sc_hd__inv_2 _20253__123 (.A(clknet_1_1__leaf__03778_),
    .Y(net247));
 sky130_fd_sc_hd__inv_2 _20254__124 (.A(clknet_1_1__leaf__03778_),
    .Y(net248));
 sky130_fd_sc_hd__inv_2 _20255__125 (.A(clknet_1_1__leaf__03778_),
    .Y(net249));
 sky130_fd_sc_hd__inv_2 _20256__126 (.A(clknet_1_1__leaf__03778_),
    .Y(net250));
 sky130_fd_sc_hd__inv_2 _20258__127 (.A(clknet_1_0__leaf__03779_),
    .Y(net251));
 sky130_fd_sc_hd__buf_1 _20257_ (.A(clknet_1_1__leaf__03464_),
    .X(_03779_));
 sky130_fd_sc_hd__inv_2 _20259__128 (.A(clknet_1_0__leaf__03779_),
    .Y(net252));
 sky130_fd_sc_hd__inv_2 _20260__129 (.A(clknet_1_0__leaf__03779_),
    .Y(net253));
 sky130_fd_sc_hd__inv_2 _20261__130 (.A(clknet_1_0__leaf__03779_),
    .Y(net254));
 sky130_fd_sc_hd__inv_2 _20262__131 (.A(clknet_1_0__leaf__03779_),
    .Y(net255));
 sky130_fd_sc_hd__inv_2 _20263__132 (.A(clknet_1_1__leaf__03779_),
    .Y(net256));
 sky130_fd_sc_hd__inv_2 _20264__133 (.A(clknet_1_1__leaf__03779_),
    .Y(net257));
 sky130_fd_sc_hd__inv_2 _20265__134 (.A(clknet_1_1__leaf__03779_),
    .Y(net258));
 sky130_fd_sc_hd__inv_2 _20266__135 (.A(clknet_1_1__leaf__03779_),
    .Y(net259));
 sky130_fd_sc_hd__inv_2 _20267__136 (.A(clknet_1_1__leaf__03779_),
    .Y(net260));
 sky130_fd_sc_hd__inv_2 _20269__137 (.A(clknet_1_0__leaf__03780_),
    .Y(net261));
 sky130_fd_sc_hd__buf_1 _20268_ (.A(clknet_1_1__leaf__03464_),
    .X(_03780_));
 sky130_fd_sc_hd__inv_2 _20270__138 (.A(clknet_1_0__leaf__03780_),
    .Y(net262));
 sky130_fd_sc_hd__inv_2 _20271__139 (.A(clknet_1_0__leaf__03780_),
    .Y(net263));
 sky130_fd_sc_hd__inv_2 _20272__140 (.A(clknet_1_0__leaf__03780_),
    .Y(net264));
 sky130_fd_sc_hd__inv_2 _20273__141 (.A(clknet_1_0__leaf__03780_),
    .Y(net265));
 sky130_fd_sc_hd__inv_2 _20274__142 (.A(clknet_1_0__leaf__03780_),
    .Y(net266));
 sky130_fd_sc_hd__inv_2 _20275__143 (.A(clknet_1_1__leaf__03780_),
    .Y(net267));
 sky130_fd_sc_hd__inv_2 _20276__144 (.A(clknet_1_1__leaf__03780_),
    .Y(net268));
 sky130_fd_sc_hd__inv_2 _20277__145 (.A(clknet_1_1__leaf__03780_),
    .Y(net269));
 sky130_fd_sc_hd__inv_2 _20278__146 (.A(clknet_1_1__leaf__03780_),
    .Y(net270));
 sky130_fd_sc_hd__inv_2 _20280__147 (.A(clknet_1_1__leaf__03781_),
    .Y(net271));
 sky130_fd_sc_hd__buf_1 _20279_ (.A(clknet_1_1__leaf__03464_),
    .X(_03781_));
 sky130_fd_sc_hd__inv_2 _20281__148 (.A(clknet_1_1__leaf__03781_),
    .Y(net272));
 sky130_fd_sc_hd__inv_2 _20282__149 (.A(clknet_1_1__leaf__03781_),
    .Y(net273));
 sky130_fd_sc_hd__inv_2 _20283__150 (.A(clknet_1_1__leaf__03781_),
    .Y(net274));
 sky130_fd_sc_hd__inv_2 _20284__151 (.A(clknet_1_1__leaf__03781_),
    .Y(net275));
 sky130_fd_sc_hd__inv_2 _20285__152 (.A(clknet_1_1__leaf__03781_),
    .Y(net276));
 sky130_fd_sc_hd__inv_2 _20286__153 (.A(clknet_1_0__leaf__03781_),
    .Y(net277));
 sky130_fd_sc_hd__inv_2 _20287__154 (.A(clknet_1_0__leaf__03781_),
    .Y(net278));
 sky130_fd_sc_hd__inv_2 _20288__155 (.A(clknet_1_0__leaf__03781_),
    .Y(net279));
 sky130_fd_sc_hd__inv_2 _20289__156 (.A(clknet_1_0__leaf__03781_),
    .Y(net280));
 sky130_fd_sc_hd__inv_2 _20291__157 (.A(clknet_1_0__leaf__03782_),
    .Y(net281));
 sky130_fd_sc_hd__buf_1 _20290_ (.A(clknet_1_1__leaf__03464_),
    .X(_03782_));
 sky130_fd_sc_hd__inv_2 _20292__158 (.A(clknet_1_0__leaf__03782_),
    .Y(net282));
 sky130_fd_sc_hd__inv_2 _20293__159 (.A(clknet_1_0__leaf__03782_),
    .Y(net283));
 sky130_fd_sc_hd__inv_2 _20294__160 (.A(clknet_1_0__leaf__03782_),
    .Y(net284));
 sky130_fd_sc_hd__inv_2 _20295__161 (.A(clknet_1_0__leaf__03782_),
    .Y(net285));
 sky130_fd_sc_hd__inv_2 _20296__162 (.A(clknet_1_1__leaf__03782_),
    .Y(net286));
 sky130_fd_sc_hd__inv_2 _20297__163 (.A(clknet_1_1__leaf__03782_),
    .Y(net287));
 sky130_fd_sc_hd__inv_2 _20298__164 (.A(clknet_1_1__leaf__03782_),
    .Y(net288));
 sky130_fd_sc_hd__inv_2 _20299__165 (.A(clknet_1_1__leaf__03782_),
    .Y(net289));
 sky130_fd_sc_hd__inv_2 _20300__166 (.A(clknet_1_1__leaf__03782_),
    .Y(net290));
 sky130_fd_sc_hd__inv_2 _20302__167 (.A(clknet_1_0__leaf__03783_),
    .Y(net291));
 sky130_fd_sc_hd__buf_1 _20301_ (.A(clknet_1_1__leaf__03464_),
    .X(_03783_));
 sky130_fd_sc_hd__inv_2 _20303__168 (.A(clknet_1_0__leaf__03783_),
    .Y(net292));
 sky130_fd_sc_hd__inv_2 _20304__169 (.A(clknet_1_0__leaf__03783_),
    .Y(net293));
 sky130_fd_sc_hd__inv_2 _20305__170 (.A(clknet_1_0__leaf__03783_),
    .Y(net294));
 sky130_fd_sc_hd__inv_2 _20306__171 (.A(clknet_1_1__leaf__03783_),
    .Y(net295));
 sky130_fd_sc_hd__inv_2 _20307__172 (.A(clknet_1_1__leaf__03783_),
    .Y(net296));
 sky130_fd_sc_hd__inv_2 _20308__173 (.A(clknet_1_1__leaf__03783_),
    .Y(net297));
 sky130_fd_sc_hd__inv_2 _20309__174 (.A(clknet_1_1__leaf__03783_),
    .Y(net298));
 sky130_fd_sc_hd__inv_2 _20310__175 (.A(clknet_1_1__leaf__03783_),
    .Y(net299));
 sky130_fd_sc_hd__inv_2 _20311__176 (.A(clknet_1_1__leaf__03783_),
    .Y(net300));
 sky130_fd_sc_hd__inv_2 _20313__177 (.A(clknet_1_0__leaf__03784_),
    .Y(net301));
 sky130_fd_sc_hd__buf_1 _20312_ (.A(clknet_1_1__leaf__03464_),
    .X(_03784_));
 sky130_fd_sc_hd__inv_2 _20314__178 (.A(clknet_1_0__leaf__03784_),
    .Y(net302));
 sky130_fd_sc_hd__inv_2 _20315__179 (.A(clknet_1_0__leaf__03784_),
    .Y(net303));
 sky130_fd_sc_hd__inv_2 _20316__180 (.A(clknet_1_0__leaf__03784_),
    .Y(net304));
 sky130_fd_sc_hd__inv_2 _20317__181 (.A(clknet_1_0__leaf__03784_),
    .Y(net305));
 sky130_fd_sc_hd__inv_2 _20318__182 (.A(clknet_1_1__leaf__03784_),
    .Y(net306));
 sky130_fd_sc_hd__inv_2 _20319__183 (.A(clknet_1_1__leaf__03784_),
    .Y(net307));
 sky130_fd_sc_hd__inv_2 _20320__184 (.A(clknet_1_1__leaf__03784_),
    .Y(net308));
 sky130_fd_sc_hd__inv_2 _20321__185 (.A(clknet_1_1__leaf__03784_),
    .Y(net309));
 sky130_fd_sc_hd__inv_2 _20322__186 (.A(clknet_1_1__leaf__03784_),
    .Y(net310));
 sky130_fd_sc_hd__inv_2 _20325__187 (.A(clknet_1_1__leaf__03786_),
    .Y(net311));
 sky130_fd_sc_hd__buf_1 _20323_ (.A(clknet_1_1__leaf__04634_),
    .X(_03785_));
 sky130_fd_sc_hd__buf_1 _20324_ (.A(clknet_1_1__leaf__03785_),
    .X(_03786_));
 sky130_fd_sc_hd__inv_2 _20326__188 (.A(clknet_1_1__leaf__03786_),
    .Y(net312));
 sky130_fd_sc_hd__inv_2 _20327__189 (.A(clknet_1_1__leaf__03786_),
    .Y(net313));
 sky130_fd_sc_hd__inv_2 _20328__190 (.A(clknet_1_1__leaf__03786_),
    .Y(net314));
 sky130_fd_sc_hd__inv_2 _20329__191 (.A(clknet_1_1__leaf__03786_),
    .Y(net315));
 sky130_fd_sc_hd__inv_2 _20330__192 (.A(clknet_1_1__leaf__03786_),
    .Y(net316));
 sky130_fd_sc_hd__inv_2 _20331__193 (.A(clknet_1_0__leaf__03786_),
    .Y(net317));
 sky130_fd_sc_hd__inv_2 _20332__194 (.A(clknet_1_0__leaf__03786_),
    .Y(net318));
 sky130_fd_sc_hd__inv_2 _20333__195 (.A(clknet_1_0__leaf__03786_),
    .Y(net319));
 sky130_fd_sc_hd__inv_2 _20334__196 (.A(clknet_1_0__leaf__03786_),
    .Y(net320));
 sky130_fd_sc_hd__inv_2 _20336__197 (.A(clknet_1_1__leaf__03787_),
    .Y(net321));
 sky130_fd_sc_hd__buf_1 _20335_ (.A(clknet_1_1__leaf__03785_),
    .X(_03787_));
 sky130_fd_sc_hd__inv_2 _20337__198 (.A(clknet_1_1__leaf__03787_),
    .Y(net322));
 sky130_fd_sc_hd__inv_2 _20338__199 (.A(clknet_1_1__leaf__03787_),
    .Y(net323));
 sky130_fd_sc_hd__inv_2 _20339__200 (.A(clknet_1_1__leaf__03787_),
    .Y(net324));
 sky130_fd_sc_hd__inv_2 _20340__201 (.A(clknet_1_1__leaf__03787_),
    .Y(net325));
 sky130_fd_sc_hd__inv_2 _20341__202 (.A(clknet_1_1__leaf__03787_),
    .Y(net326));
 sky130_fd_sc_hd__inv_2 _20342__203 (.A(clknet_1_0__leaf__03787_),
    .Y(net327));
 sky130_fd_sc_hd__inv_2 _20343__204 (.A(clknet_1_0__leaf__03787_),
    .Y(net328));
 sky130_fd_sc_hd__inv_2 _20344__205 (.A(clknet_1_0__leaf__03787_),
    .Y(net329));
 sky130_fd_sc_hd__inv_2 _20345__206 (.A(clknet_1_0__leaf__03787_),
    .Y(net330));
 sky130_fd_sc_hd__inv_2 _20347__207 (.A(clknet_1_0__leaf__03788_),
    .Y(net331));
 sky130_fd_sc_hd__buf_1 _20346_ (.A(clknet_1_1__leaf__03785_),
    .X(_03788_));
 sky130_fd_sc_hd__inv_2 _20348__208 (.A(clknet_1_0__leaf__03788_),
    .Y(net332));
 sky130_fd_sc_hd__inv_2 _20349__209 (.A(clknet_1_0__leaf__03788_),
    .Y(net333));
 sky130_fd_sc_hd__inv_2 _20350__210 (.A(clknet_1_0__leaf__03788_),
    .Y(net334));
 sky130_fd_sc_hd__inv_2 _20351__211 (.A(clknet_1_0__leaf__03788_),
    .Y(net335));
 sky130_fd_sc_hd__inv_2 _20352__212 (.A(clknet_1_1__leaf__03788_),
    .Y(net336));
 sky130_fd_sc_hd__inv_2 _20353__213 (.A(clknet_1_1__leaf__03788_),
    .Y(net337));
 sky130_fd_sc_hd__inv_2 _20354__214 (.A(clknet_1_1__leaf__03788_),
    .Y(net338));
 sky130_fd_sc_hd__inv_2 _20355__215 (.A(clknet_1_1__leaf__03788_),
    .Y(net339));
 sky130_fd_sc_hd__inv_2 _20356__216 (.A(clknet_1_1__leaf__03788_),
    .Y(net340));
 sky130_fd_sc_hd__inv_2 _20358__217 (.A(clknet_1_0__leaf__03789_),
    .Y(net341));
 sky130_fd_sc_hd__buf_1 _20357_ (.A(clknet_1_1__leaf__03785_),
    .X(_03789_));
 sky130_fd_sc_hd__inv_2 _20359__218 (.A(clknet_1_0__leaf__03789_),
    .Y(net342));
 sky130_fd_sc_hd__inv_2 _20360__219 (.A(clknet_1_1__leaf__03789_),
    .Y(net343));
 sky130_fd_sc_hd__inv_2 _20361__220 (.A(clknet_1_0__leaf__03789_),
    .Y(net344));
 sky130_fd_sc_hd__inv_2 _20362__221 (.A(clknet_1_0__leaf__03789_),
    .Y(net345));
 sky130_fd_sc_hd__inv_2 _20363__222 (.A(clknet_1_0__leaf__03789_),
    .Y(net346));
 sky130_fd_sc_hd__inv_2 _20364__223 (.A(clknet_1_0__leaf__03789_),
    .Y(net347));
 sky130_fd_sc_hd__inv_2 _20365__224 (.A(clknet_1_1__leaf__03789_),
    .Y(net348));
 sky130_fd_sc_hd__inv_2 _20366__225 (.A(clknet_1_1__leaf__03789_),
    .Y(net349));
 sky130_fd_sc_hd__inv_2 _20367__226 (.A(clknet_1_1__leaf__03789_),
    .Y(net350));
 sky130_fd_sc_hd__inv_2 _20369__227 (.A(clknet_1_0__leaf__03790_),
    .Y(net351));
 sky130_fd_sc_hd__buf_1 _20368_ (.A(clknet_1_0__leaf__03785_),
    .X(_03790_));
 sky130_fd_sc_hd__inv_2 _20370__228 (.A(clknet_1_0__leaf__03790_),
    .Y(net352));
 sky130_fd_sc_hd__inv_2 _20371__229 (.A(clknet_1_0__leaf__03790_),
    .Y(net353));
 sky130_fd_sc_hd__inv_2 _20372__230 (.A(clknet_1_0__leaf__03790_),
    .Y(net354));
 sky130_fd_sc_hd__inv_2 _20373__231 (.A(clknet_1_0__leaf__03790_),
    .Y(net355));
 sky130_fd_sc_hd__inv_2 _20374__232 (.A(clknet_1_0__leaf__03790_),
    .Y(net356));
 sky130_fd_sc_hd__inv_2 _20375__233 (.A(clknet_1_1__leaf__03790_),
    .Y(net357));
 sky130_fd_sc_hd__inv_2 _20376__234 (.A(clknet_1_1__leaf__03790_),
    .Y(net358));
 sky130_fd_sc_hd__inv_2 _20377__235 (.A(clknet_1_1__leaf__03790_),
    .Y(net359));
 sky130_fd_sc_hd__inv_2 _20378__236 (.A(clknet_1_1__leaf__03790_),
    .Y(net360));
 sky130_fd_sc_hd__inv_2 _20380__237 (.A(clknet_1_1__leaf__03791_),
    .Y(net361));
 sky130_fd_sc_hd__buf_1 _20379_ (.A(clknet_1_0__leaf__03785_),
    .X(_03791_));
 sky130_fd_sc_hd__inv_2 _20381__238 (.A(clknet_1_1__leaf__03791_),
    .Y(net362));
 sky130_fd_sc_hd__inv_2 _20382__239 (.A(clknet_1_1__leaf__03791_),
    .Y(net363));
 sky130_fd_sc_hd__inv_2 _20383__240 (.A(clknet_1_1__leaf__03791_),
    .Y(net364));
 sky130_fd_sc_hd__inv_2 _20384__241 (.A(clknet_1_1__leaf__03791_),
    .Y(net365));
 sky130_fd_sc_hd__inv_2 _20385__242 (.A(clknet_1_1__leaf__03791_),
    .Y(net366));
 sky130_fd_sc_hd__inv_2 _20386__243 (.A(clknet_1_0__leaf__03791_),
    .Y(net367));
 sky130_fd_sc_hd__inv_2 _20387__244 (.A(clknet_1_0__leaf__03791_),
    .Y(net368));
 sky130_fd_sc_hd__inv_2 _20388__245 (.A(clknet_1_0__leaf__03791_),
    .Y(net369));
 sky130_fd_sc_hd__inv_2 _20389__246 (.A(clknet_1_0__leaf__03791_),
    .Y(net370));
 sky130_fd_sc_hd__inv_2 _20391__247 (.A(clknet_1_1__leaf__03792_),
    .Y(net371));
 sky130_fd_sc_hd__buf_1 _20390_ (.A(clknet_1_0__leaf__03785_),
    .X(_03792_));
 sky130_fd_sc_hd__inv_2 _20392__248 (.A(clknet_1_1__leaf__03792_),
    .Y(net372));
 sky130_fd_sc_hd__inv_2 _20393__249 (.A(clknet_1_1__leaf__03792_),
    .Y(net373));
 sky130_fd_sc_hd__inv_2 _20394__250 (.A(clknet_1_1__leaf__03792_),
    .Y(net374));
 sky130_fd_sc_hd__inv_2 _20395__251 (.A(clknet_1_1__leaf__03792_),
    .Y(net375));
 sky130_fd_sc_hd__inv_2 _20396__252 (.A(clknet_1_0__leaf__03792_),
    .Y(net376));
 sky130_fd_sc_hd__inv_2 _20397__253 (.A(clknet_1_0__leaf__03792_),
    .Y(net377));
 sky130_fd_sc_hd__inv_2 _20398__254 (.A(clknet_1_0__leaf__03792_),
    .Y(net378));
 sky130_fd_sc_hd__inv_2 _20399__255 (.A(clknet_1_0__leaf__03792_),
    .Y(net379));
 sky130_fd_sc_hd__inv_2 _20400__256 (.A(clknet_1_0__leaf__03792_),
    .Y(net380));
 sky130_fd_sc_hd__inv_2 _20402__257 (.A(clknet_1_0__leaf__03793_),
    .Y(net381));
 sky130_fd_sc_hd__buf_1 _20401_ (.A(clknet_1_0__leaf__03785_),
    .X(_03793_));
 sky130_fd_sc_hd__inv_2 _20403__258 (.A(clknet_1_0__leaf__03793_),
    .Y(net382));
 sky130_fd_sc_hd__inv_2 _20404__259 (.A(clknet_1_0__leaf__03793_),
    .Y(net383));
 sky130_fd_sc_hd__inv_2 _20405__260 (.A(clknet_1_0__leaf__03793_),
    .Y(net384));
 sky130_fd_sc_hd__inv_2 _20406__261 (.A(clknet_1_0__leaf__03793_),
    .Y(net385));
 sky130_fd_sc_hd__inv_2 _20407__262 (.A(clknet_1_0__leaf__03793_),
    .Y(net386));
 sky130_fd_sc_hd__inv_2 _20408__263 (.A(clknet_1_1__leaf__03793_),
    .Y(net387));
 sky130_fd_sc_hd__inv_2 _20409__264 (.A(clknet_1_1__leaf__03793_),
    .Y(net388));
 sky130_fd_sc_hd__inv_2 _20410__265 (.A(clknet_1_1__leaf__03793_),
    .Y(net389));
 sky130_fd_sc_hd__inv_2 _20411__266 (.A(clknet_1_1__leaf__03793_),
    .Y(net390));
 sky130_fd_sc_hd__inv_2 _20413__267 (.A(clknet_1_1__leaf__03794_),
    .Y(net391));
 sky130_fd_sc_hd__buf_1 _20412_ (.A(clknet_1_0__leaf__03785_),
    .X(_03794_));
 sky130_fd_sc_hd__inv_2 _20414__268 (.A(clknet_1_1__leaf__03794_),
    .Y(net392));
 sky130_fd_sc_hd__inv_2 _20415__269 (.A(clknet_1_1__leaf__03794_),
    .Y(net393));
 sky130_fd_sc_hd__inv_2 _20416__270 (.A(clknet_1_1__leaf__03794_),
    .Y(net394));
 sky130_fd_sc_hd__inv_2 _20417__271 (.A(clknet_1_1__leaf__03794_),
    .Y(net395));
 sky130_fd_sc_hd__inv_2 _20418__272 (.A(clknet_1_1__leaf__03794_),
    .Y(net396));
 sky130_fd_sc_hd__inv_2 _20419__273 (.A(clknet_1_0__leaf__03794_),
    .Y(net397));
 sky130_fd_sc_hd__inv_2 _20420__274 (.A(clknet_1_0__leaf__03794_),
    .Y(net398));
 sky130_fd_sc_hd__inv_2 _20421__275 (.A(clknet_1_0__leaf__03794_),
    .Y(net399));
 sky130_fd_sc_hd__inv_2 _20422__276 (.A(clknet_1_0__leaf__03794_),
    .Y(net400));
 sky130_fd_sc_hd__inv_2 _20424__277 (.A(clknet_1_1__leaf__03795_),
    .Y(net401));
 sky130_fd_sc_hd__buf_1 _20423_ (.A(clknet_1_0__leaf__03785_),
    .X(_03795_));
 sky130_fd_sc_hd__inv_2 _20425__278 (.A(clknet_1_0__leaf__03795_),
    .Y(net402));
 sky130_fd_sc_hd__inv_2 _20426__279 (.A(clknet_1_0__leaf__03795_),
    .Y(net403));
 sky130_fd_sc_hd__inv_2 _20427__280 (.A(clknet_1_0__leaf__03795_),
    .Y(net404));
 sky130_fd_sc_hd__inv_2 _20428__281 (.A(clknet_1_0__leaf__03795_),
    .Y(net405));
 sky130_fd_sc_hd__inv_2 _20429__282 (.A(clknet_1_0__leaf__03795_),
    .Y(net406));
 sky130_fd_sc_hd__inv_2 _20430__283 (.A(clknet_1_1__leaf__03795_),
    .Y(net407));
 sky130_fd_sc_hd__inv_2 _20431__284 (.A(clknet_1_1__leaf__03795_),
    .Y(net408));
 sky130_fd_sc_hd__inv_2 _20432__285 (.A(clknet_1_1__leaf__03795_),
    .Y(net409));
 sky130_fd_sc_hd__inv_2 _20433__286 (.A(clknet_1_1__leaf__03795_),
    .Y(net410));
 sky130_fd_sc_hd__inv_2 _20436__287 (.A(clknet_1_0__leaf__03797_),
    .Y(net411));
 sky130_fd_sc_hd__buf_1 _20434_ (.A(clknet_1_1__leaf__04634_),
    .X(_03796_));
 sky130_fd_sc_hd__buf_1 _20435_ (.A(clknet_1_1__leaf__03796_),
    .X(_03797_));
 sky130_fd_sc_hd__inv_2 _20437__288 (.A(clknet_1_0__leaf__03797_),
    .Y(net412));
 sky130_fd_sc_hd__inv_2 _20438__289 (.A(clknet_1_0__leaf__03797_),
    .Y(net413));
 sky130_fd_sc_hd__inv_2 _20439__290 (.A(clknet_1_0__leaf__03797_),
    .Y(net414));
 sky130_fd_sc_hd__inv_2 _20440__291 (.A(clknet_1_1__leaf__03797_),
    .Y(net415));
 sky130_fd_sc_hd__inv_2 _20441__292 (.A(clknet_1_1__leaf__03797_),
    .Y(net416));
 sky130_fd_sc_hd__inv_2 _20442__293 (.A(clknet_1_1__leaf__03797_),
    .Y(net417));
 sky130_fd_sc_hd__inv_2 _20443__294 (.A(clknet_1_1__leaf__03797_),
    .Y(net418));
 sky130_fd_sc_hd__inv_2 _20444__295 (.A(clknet_1_1__leaf__03797_),
    .Y(net419));
 sky130_fd_sc_hd__inv_2 _20445__296 (.A(clknet_1_1__leaf__03797_),
    .Y(net420));
 sky130_fd_sc_hd__inv_2 _20447__297 (.A(clknet_1_1__leaf__03798_),
    .Y(net421));
 sky130_fd_sc_hd__buf_1 _20446_ (.A(clknet_1_1__leaf__03796_),
    .X(_03798_));
 sky130_fd_sc_hd__inv_2 _20448__298 (.A(clknet_1_1__leaf__03798_),
    .Y(net422));
 sky130_fd_sc_hd__inv_2 _20449__299 (.A(clknet_1_1__leaf__03798_),
    .Y(net423));
 sky130_fd_sc_hd__inv_2 _20450__300 (.A(clknet_1_1__leaf__03798_),
    .Y(net424));
 sky130_fd_sc_hd__inv_2 _20451__301 (.A(clknet_1_1__leaf__03798_),
    .Y(net425));
 sky130_fd_sc_hd__inv_2 _20452__302 (.A(clknet_1_1__leaf__03798_),
    .Y(net426));
 sky130_fd_sc_hd__inv_2 _20453__303 (.A(clknet_1_0__leaf__03798_),
    .Y(net427));
 sky130_fd_sc_hd__inv_2 _20454__304 (.A(clknet_1_0__leaf__03798_),
    .Y(net428));
 sky130_fd_sc_hd__inv_2 _20455__305 (.A(clknet_1_0__leaf__03798_),
    .Y(net429));
 sky130_fd_sc_hd__inv_2 _20456__306 (.A(clknet_1_0__leaf__03798_),
    .Y(net430));
 sky130_fd_sc_hd__inv_2 _20458__307 (.A(clknet_1_1__leaf__03799_),
    .Y(net431));
 sky130_fd_sc_hd__buf_1 _20457_ (.A(clknet_1_1__leaf__03796_),
    .X(_03799_));
 sky130_fd_sc_hd__inv_2 _20459__308 (.A(clknet_1_1__leaf__03799_),
    .Y(net432));
 sky130_fd_sc_hd__inv_2 _20460__309 (.A(clknet_1_1__leaf__03799_),
    .Y(net433));
 sky130_fd_sc_hd__inv_2 _20461__310 (.A(clknet_1_1__leaf__03799_),
    .Y(net434));
 sky130_fd_sc_hd__inv_2 _20462__311 (.A(clknet_1_1__leaf__03799_),
    .Y(net435));
 sky130_fd_sc_hd__inv_2 _20463__312 (.A(clknet_1_0__leaf__03799_),
    .Y(net436));
 sky130_fd_sc_hd__inv_2 _20464__313 (.A(clknet_1_0__leaf__03799_),
    .Y(net437));
 sky130_fd_sc_hd__inv_2 _20465__314 (.A(clknet_1_0__leaf__03799_),
    .Y(net438));
 sky130_fd_sc_hd__inv_2 _20466__315 (.A(clknet_1_0__leaf__03799_),
    .Y(net439));
 sky130_fd_sc_hd__inv_2 _20467__316 (.A(clknet_1_0__leaf__03799_),
    .Y(net440));
 sky130_fd_sc_hd__inv_2 _20469__317 (.A(clknet_1_0__leaf__03800_),
    .Y(net441));
 sky130_fd_sc_hd__buf_1 _20468_ (.A(clknet_1_1__leaf__03796_),
    .X(_03800_));
 sky130_fd_sc_hd__inv_2 _20470__318 (.A(clknet_1_0__leaf__03800_),
    .Y(net442));
 sky130_fd_sc_hd__inv_2 _20471__319 (.A(clknet_1_0__leaf__03800_),
    .Y(net443));
 sky130_fd_sc_hd__inv_2 _20472__320 (.A(clknet_1_0__leaf__03800_),
    .Y(net444));
 sky130_fd_sc_hd__inv_2 _20473__321 (.A(clknet_1_0__leaf__03800_),
    .Y(net445));
 sky130_fd_sc_hd__inv_2 _20474__322 (.A(clknet_1_0__leaf__03800_),
    .Y(net446));
 sky130_fd_sc_hd__inv_2 _20475__323 (.A(clknet_1_1__leaf__03800_),
    .Y(net447));
 sky130_fd_sc_hd__inv_2 _20476__324 (.A(clknet_1_1__leaf__03800_),
    .Y(net448));
 sky130_fd_sc_hd__inv_2 _20477__325 (.A(clknet_1_1__leaf__03800_),
    .Y(net449));
 sky130_fd_sc_hd__inv_2 _20478__326 (.A(clknet_1_1__leaf__03800_),
    .Y(net450));
 sky130_fd_sc_hd__inv_2 _20480__327 (.A(clknet_1_1__leaf__03801_),
    .Y(net451));
 sky130_fd_sc_hd__buf_1 _20479_ (.A(clknet_1_1__leaf__03796_),
    .X(_03801_));
 sky130_fd_sc_hd__inv_2 _20481__328 (.A(clknet_1_1__leaf__03801_),
    .Y(net452));
 sky130_fd_sc_hd__inv_2 _20482__329 (.A(clknet_1_0__leaf__03801_),
    .Y(net453));
 sky130_fd_sc_hd__inv_2 _20483__330 (.A(clknet_1_0__leaf__03801_),
    .Y(net454));
 sky130_fd_sc_hd__inv_2 _20484__331 (.A(clknet_1_0__leaf__03801_),
    .Y(net455));
 sky130_fd_sc_hd__inv_2 _20485__332 (.A(clknet_1_0__leaf__03801_),
    .Y(net456));
 sky130_fd_sc_hd__inv_2 _20486__333 (.A(clknet_1_0__leaf__03801_),
    .Y(net457));
 sky130_fd_sc_hd__inv_2 _20487__334 (.A(clknet_1_1__leaf__03801_),
    .Y(net458));
 sky130_fd_sc_hd__inv_2 _20488__335 (.A(clknet_1_1__leaf__03801_),
    .Y(net459));
 sky130_fd_sc_hd__inv_2 _20489__336 (.A(clknet_1_1__leaf__03801_),
    .Y(net460));
 sky130_fd_sc_hd__inv_2 _20491__337 (.A(clknet_1_0__leaf__03802_),
    .Y(net461));
 sky130_fd_sc_hd__buf_1 _20490_ (.A(clknet_1_1__leaf__03796_),
    .X(_03802_));
 sky130_fd_sc_hd__inv_2 _20492__338 (.A(clknet_1_0__leaf__03802_),
    .Y(net462));
 sky130_fd_sc_hd__inv_2 _20493__339 (.A(clknet_1_0__leaf__03802_),
    .Y(net463));
 sky130_fd_sc_hd__inv_2 _20494__340 (.A(clknet_1_1__leaf__03802_),
    .Y(net464));
 sky130_fd_sc_hd__inv_2 _20495__341 (.A(clknet_1_1__leaf__03802_),
    .Y(net465));
 sky130_fd_sc_hd__inv_2 _20496__342 (.A(clknet_1_1__leaf__03802_),
    .Y(net466));
 sky130_fd_sc_hd__inv_2 _20497__343 (.A(clknet_1_1__leaf__03802_),
    .Y(net467));
 sky130_fd_sc_hd__inv_2 _20498__344 (.A(clknet_1_0__leaf__03802_),
    .Y(net468));
 sky130_fd_sc_hd__inv_2 _20499__345 (.A(clknet_1_0__leaf__03802_),
    .Y(net469));
 sky130_fd_sc_hd__inv_2 _20500__346 (.A(clknet_1_0__leaf__03802_),
    .Y(net470));
 sky130_fd_sc_hd__inv_2 _20502__347 (.A(clknet_1_0__leaf__03803_),
    .Y(net471));
 sky130_fd_sc_hd__buf_1 _20501_ (.A(clknet_1_0__leaf__03796_),
    .X(_03803_));
 sky130_fd_sc_hd__inv_2 _20503__348 (.A(clknet_1_0__leaf__03803_),
    .Y(net472));
 sky130_fd_sc_hd__inv_2 _20504__349 (.A(clknet_1_0__leaf__03803_),
    .Y(net473));
 sky130_fd_sc_hd__inv_2 _20505__350 (.A(clknet_1_0__leaf__03803_),
    .Y(net474));
 sky130_fd_sc_hd__inv_2 _20506__351 (.A(clknet_1_0__leaf__03803_),
    .Y(net475));
 sky130_fd_sc_hd__inv_2 _20507__352 (.A(clknet_1_1__leaf__03803_),
    .Y(net476));
 sky130_fd_sc_hd__inv_2 _20508__353 (.A(clknet_1_1__leaf__03803_),
    .Y(net477));
 sky130_fd_sc_hd__inv_2 _20509__354 (.A(clknet_1_1__leaf__03803_),
    .Y(net478));
 sky130_fd_sc_hd__inv_2 _20510__355 (.A(clknet_1_1__leaf__03803_),
    .Y(net479));
 sky130_fd_sc_hd__inv_2 _20511__356 (.A(clknet_1_1__leaf__03803_),
    .Y(net480));
 sky130_fd_sc_hd__inv_2 _20513__357 (.A(clknet_1_0__leaf__03804_),
    .Y(net481));
 sky130_fd_sc_hd__buf_1 _20512_ (.A(clknet_1_0__leaf__03796_),
    .X(_03804_));
 sky130_fd_sc_hd__inv_2 _20514__358 (.A(clknet_1_1__leaf__03804_),
    .Y(net482));
 sky130_fd_sc_hd__inv_2 _20515__359 (.A(clknet_1_1__leaf__03804_),
    .Y(net483));
 sky130_fd_sc_hd__inv_2 _20516__360 (.A(clknet_1_1__leaf__03804_),
    .Y(net484));
 sky130_fd_sc_hd__inv_2 _20517__361 (.A(clknet_1_1__leaf__03804_),
    .Y(net485));
 sky130_fd_sc_hd__inv_2 _20518__362 (.A(clknet_1_1__leaf__03804_),
    .Y(net486));
 sky130_fd_sc_hd__inv_2 _20519__363 (.A(clknet_1_0__leaf__03804_),
    .Y(net487));
 sky130_fd_sc_hd__inv_2 _20520__364 (.A(clknet_1_0__leaf__03804_),
    .Y(net488));
 sky130_fd_sc_hd__inv_2 _20521__365 (.A(clknet_1_0__leaf__03804_),
    .Y(net489));
 sky130_fd_sc_hd__inv_2 _20522__366 (.A(clknet_1_0__leaf__03804_),
    .Y(net490));
 sky130_fd_sc_hd__inv_2 _20524__367 (.A(clknet_1_1__leaf__03805_),
    .Y(net491));
 sky130_fd_sc_hd__buf_1 _20523_ (.A(clknet_1_0__leaf__03796_),
    .X(_03805_));
 sky130_fd_sc_hd__inv_2 _20525__368 (.A(clknet_1_1__leaf__03805_),
    .Y(net492));
 sky130_fd_sc_hd__inv_2 _20526__369 (.A(clknet_1_1__leaf__03805_),
    .Y(net493));
 sky130_fd_sc_hd__inv_2 _20527__370 (.A(clknet_1_1__leaf__03805_),
    .Y(net494));
 sky130_fd_sc_hd__inv_2 _20528__371 (.A(clknet_1_0__leaf__03805_),
    .Y(net495));
 sky130_fd_sc_hd__inv_2 _20529__372 (.A(clknet_1_1__leaf__03805_),
    .Y(net496));
 sky130_fd_sc_hd__inv_2 _20530__373 (.A(clknet_1_0__leaf__03805_),
    .Y(net497));
 sky130_fd_sc_hd__inv_2 _20531__374 (.A(clknet_1_0__leaf__03805_),
    .Y(net498));
 sky130_fd_sc_hd__inv_2 _20532__375 (.A(clknet_1_0__leaf__03805_),
    .Y(net499));
 sky130_fd_sc_hd__inv_2 _20533__376 (.A(clknet_1_0__leaf__03805_),
    .Y(net500));
 sky130_fd_sc_hd__inv_2 _20535__377 (.A(clknet_1_1__leaf__03806_),
    .Y(net501));
 sky130_fd_sc_hd__buf_1 _20534_ (.A(clknet_1_0__leaf__03796_),
    .X(_03806_));
 sky130_fd_sc_hd__inv_2 _20536__378 (.A(clknet_1_1__leaf__03806_),
    .Y(net502));
 sky130_fd_sc_hd__inv_2 _20537__379 (.A(clknet_1_1__leaf__03806_),
    .Y(net503));
 sky130_fd_sc_hd__inv_2 _20538__380 (.A(clknet_1_1__leaf__03806_),
    .Y(net504));
 sky130_fd_sc_hd__inv_2 _20539__381 (.A(clknet_1_1__leaf__03806_),
    .Y(net505));
 sky130_fd_sc_hd__inv_2 _20540__382 (.A(clknet_1_1__leaf__03806_),
    .Y(net506));
 sky130_fd_sc_hd__inv_2 _20541__383 (.A(clknet_1_0__leaf__03806_),
    .Y(net507));
 sky130_fd_sc_hd__inv_2 _20542__384 (.A(clknet_1_0__leaf__03806_),
    .Y(net508));
 sky130_fd_sc_hd__inv_2 _20543__385 (.A(clknet_1_0__leaf__03806_),
    .Y(net509));
 sky130_fd_sc_hd__inv_2 _20544__386 (.A(clknet_1_0__leaf__03806_),
    .Y(net510));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__buf_1 _20545_ (.A(clknet_1_0__leaf__04634_),
    .X(_03807_));
 sky130_fd_sc_hd__inv_2 _20547__8 (.A(clknet_1_1__leaf__03807_),
    .Y(net132));
 sky130_fd_sc_hd__inv_2 _20548__9 (.A(clknet_1_1__leaf__03807_),
    .Y(net133));
 sky130_fd_sc_hd__inv_2 _20549__10 (.A(clknet_1_1__leaf__03807_),
    .Y(net134));
 sky130_fd_sc_hd__inv_2 _20550__11 (.A(clknet_1_1__leaf__03807_),
    .Y(net135));
 sky130_fd_sc_hd__inv_2 _20551__12 (.A(clknet_1_0__leaf__03807_),
    .Y(net136));
 sky130_fd_sc_hd__inv_2 _20552__13 (.A(clknet_1_0__leaf__03807_),
    .Y(net137));
 sky130_fd_sc_hd__inv_2 _20553__14 (.A(clknet_1_0__leaf__03807_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _20554__15 (.A(clknet_1_0__leaf__03807_),
    .Y(net139));
 sky130_fd_sc_hd__inv_2 _20555__16 (.A(clknet_1_0__leaf__03807_),
    .Y(net140));
 sky130_fd_sc_hd__inv_2 _20557__17 (.A(clknet_1_0__leaf__03808_),
    .Y(net141));
 sky130_fd_sc_hd__buf_1 _20556_ (.A(clknet_1_1__leaf__04634_),
    .X(_03808_));
 sky130_fd_sc_hd__inv_2 _20558__18 (.A(clknet_1_0__leaf__03808_),
    .Y(net142));
 sky130_fd_sc_hd__inv_2 _20559__19 (.A(clknet_1_1__leaf__03808_),
    .Y(net143));
 sky130_fd_sc_hd__inv_2 _20560__20 (.A(clknet_1_1__leaf__03808_),
    .Y(net144));
 sky130_fd_sc_hd__inv_2 _20561__21 (.A(clknet_1_1__leaf__03808_),
    .Y(net145));
 sky130_fd_sc_hd__inv_2 _20562__22 (.A(clknet_1_1__leaf__03808_),
    .Y(net146));
 sky130_fd_sc_hd__inv_2 _20563__23 (.A(clknet_1_0__leaf__03808_),
    .Y(net147));
 sky130_fd_sc_hd__inv_2 _20564__24 (.A(clknet_1_0__leaf__03808_),
    .Y(net148));
 sky130_fd_sc_hd__inv_2 _20565__25 (.A(clknet_1_0__leaf__03808_),
    .Y(net149));
 sky130_fd_sc_hd__inv_2 _20566__26 (.A(clknet_1_0__leaf__03808_),
    .Y(net150));
 sky130_fd_sc_hd__inv_2 _19645__27 (.A(clknet_1_1__leaf__03458_),
    .Y(net151));
 sky130_fd_sc_hd__inv_2 _20568__4 (.A(clknet_1_1__leaf__03457_),
    .Y(net128));
 sky130_fd_sc_hd__inv_2 _20569__5 (.A(clknet_1_1__leaf__03457_),
    .Y(net129));
 sky130_fd_sc_hd__inv_2 _20570__6 (.A(clknet_1_1__leaf__03457_),
    .Y(net130));
 sky130_fd_sc_hd__inv_2 _20546__7 (.A(clknet_1_1__leaf__03807_),
    .Y(net131));
 sky130_fd_sc_hd__nor2_1 _20571_ (.A(\gpout5.clk_div[0] ),
    .B(net63),
    .Y(_01598_));
 sky130_fd_sc_hd__nand2_1 _20572_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .Y(_03809_));
 sky130_fd_sc_hd__or2_1 _20573_ (.A(\gpout5.clk_div[1] ),
    .B(\gpout5.clk_div[0] ),
    .X(_03810_));
 sky130_fd_sc_hd__and3_1 _20574_ (.A(_03728_),
    .B(_03809_),
    .C(_03810_),
    .X(_03811_));
 sky130_fd_sc_hd__clkbuf_1 _20575_ (.A(_03811_),
    .X(_01599_));
 sky130_fd_sc_hd__nand2_1 _20576_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .Y(_03812_));
 sky130_fd_sc_hd__or2_1 _20577_ (.A(\rbzero.traced_texa[-11] ),
    .B(\rbzero.texV[-11] ),
    .X(_03813_));
 sky130_fd_sc_hd__clkbuf_4 _20578_ (.A(_09734_),
    .X(_03814_));
 sky130_fd_sc_hd__a32o_1 _20579_ (.A1(_03734_),
    .A2(_03812_),
    .A3(_03813_),
    .B1(_03814_),
    .B2(\rbzero.texV[-11] ),
    .X(_01600_));
 sky130_fd_sc_hd__or2_1 _20580_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .X(_03815_));
 sky130_fd_sc_hd__nand2_1 _20581_ (.A(\rbzero.traced_texa[-10] ),
    .B(\rbzero.texV[-10] ),
    .Y(_03816_));
 sky130_fd_sc_hd__nand3b_1 _20582_ (.A_N(_03812_),
    .B(_03815_),
    .C(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__a21bo_1 _20583_ (.A1(_03815_),
    .A2(_03816_),
    .B1_N(_03812_),
    .X(_03818_));
 sky130_fd_sc_hd__a32o_1 _20584_ (.A1(_03734_),
    .A2(_03817_),
    .A3(_03818_),
    .B1(_03814_),
    .B2(\rbzero.texV[-10] ),
    .X(_01601_));
 sky130_fd_sc_hd__buf_4 _20585_ (.A(_09732_),
    .X(_03819_));
 sky130_fd_sc_hd__and2_1 _20586_ (.A(_03816_),
    .B(_03817_),
    .X(_03820_));
 sky130_fd_sc_hd__nor2_1 _20587_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_03821_));
 sky130_fd_sc_hd__nand2_1 _20588_ (.A(\rbzero.traced_texa[-9] ),
    .B(\rbzero.texV[-9] ),
    .Y(_03822_));
 sky130_fd_sc_hd__and2b_1 _20589_ (.A_N(_03821_),
    .B(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__xnor2_1 _20590_ (.A(_03820_),
    .B(_03823_),
    .Y(_03824_));
 sky130_fd_sc_hd__a22o_1 _20591_ (.A1(\rbzero.texV[-9] ),
    .A2(_03695_),
    .B1(_03819_),
    .B2(_03824_),
    .X(_01602_));
 sky130_fd_sc_hd__or2_1 _20592_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .X(_03825_));
 sky130_fd_sc_hd__nand2_1 _20593_ (.A(\rbzero.traced_texa[-8] ),
    .B(\rbzero.texV[-8] ),
    .Y(_03826_));
 sky130_fd_sc_hd__nand2_1 _20594_ (.A(_03825_),
    .B(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__o21ai_1 _20595_ (.A1(_03820_),
    .A2(_03821_),
    .B1(_03822_),
    .Y(_03828_));
 sky130_fd_sc_hd__xnor2_1 _20596_ (.A(_03827_),
    .B(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__a22o_1 _20597_ (.A1(\rbzero.texV[-8] ),
    .A2(_03695_),
    .B1(_03819_),
    .B2(_03829_),
    .X(_01603_));
 sky130_fd_sc_hd__nor2_1 _20598_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .Y(_03830_));
 sky130_fd_sc_hd__and2_1 _20599_ (.A(\rbzero.traced_texa[-7] ),
    .B(\rbzero.texV[-7] ),
    .X(_03831_));
 sky130_fd_sc_hd__a21boi_1 _20600_ (.A1(_03825_),
    .A2(_03828_),
    .B1_N(_03826_),
    .Y(_03832_));
 sky130_fd_sc_hd__o21ai_1 _20601_ (.A1(_03830_),
    .A2(_03831_),
    .B1(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__or3_1 _20602_ (.A(_03830_),
    .B(_03831_),
    .C(_03832_),
    .X(_03834_));
 sky130_fd_sc_hd__a32o_1 _20603_ (.A1(_03734_),
    .A2(_03833_),
    .A3(_03834_),
    .B1(_03814_),
    .B2(\rbzero.texV[-7] ),
    .X(_01604_));
 sky130_fd_sc_hd__xnor2_1 _20604_ (.A(\rbzero.traced_texa[-6] ),
    .B(\rbzero.texV[-6] ),
    .Y(_03835_));
 sky130_fd_sc_hd__o21bai_1 _20605_ (.A1(_03830_),
    .A2(_03832_),
    .B1_N(_03831_),
    .Y(_03836_));
 sky130_fd_sc_hd__xnor2_1 _20606_ (.A(_03835_),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__a22o_1 _20607_ (.A1(\rbzero.texV[-6] ),
    .A2(_03695_),
    .B1(_03819_),
    .B2(_03837_),
    .X(_01605_));
 sky130_fd_sc_hd__nor2_1 _20608_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .Y(_03838_));
 sky130_fd_sc_hd__nand2_1 _20609_ (.A(\rbzero.traced_texa[-5] ),
    .B(\rbzero.texV[-5] ),
    .Y(_03839_));
 sky130_fd_sc_hd__and2b_1 _20610_ (.A_N(_03838_),
    .B(_03839_),
    .X(_03840_));
 sky130_fd_sc_hd__a21o_1 _20611_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(\rbzero.texV[-6] ),
    .B1(_03836_),
    .X(_03841_));
 sky130_fd_sc_hd__o21ai_1 _20612_ (.A1(\rbzero.traced_texa[-6] ),
    .A2(\rbzero.texV[-6] ),
    .B1(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__xnor2_1 _20613_ (.A(_03840_),
    .B(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__a22o_1 _20614_ (.A1(\rbzero.texV[-5] ),
    .A2(_03814_),
    .B1(_03819_),
    .B2(_03843_),
    .X(_01606_));
 sky130_fd_sc_hd__or2_1 _20615_ (.A(\rbzero.traced_texa[-4] ),
    .B(\rbzero.texV[-4] ),
    .X(_03844_));
 sky130_fd_sc_hd__nand2_1 _20616_ (.A(\rbzero.traced_texa[-4] ),
    .B(\rbzero.texV[-4] ),
    .Y(_03845_));
 sky130_fd_sc_hd__o21ai_1 _20617_ (.A1(_03838_),
    .A2(_03842_),
    .B1(_03839_),
    .Y(_03846_));
 sky130_fd_sc_hd__nand3_1 _20618_ (.A(_03844_),
    .B(_03845_),
    .C(_03846_),
    .Y(_03847_));
 sky130_fd_sc_hd__a21o_1 _20619_ (.A1(_03844_),
    .A2(_03845_),
    .B1(_03846_),
    .X(_03848_));
 sky130_fd_sc_hd__a32o_1 _20620_ (.A1(_03734_),
    .A2(_03847_),
    .A3(_03848_),
    .B1(_03740_),
    .B2(\rbzero.texV[-4] ),
    .X(_01607_));
 sky130_fd_sc_hd__nor2_1 _20621_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_03849_));
 sky130_fd_sc_hd__nand2_1 _20622_ (.A(\rbzero.traced_texa[-3] ),
    .B(\rbzero.texV[-3] ),
    .Y(_03850_));
 sky130_fd_sc_hd__and2b_1 _20623_ (.A_N(_03849_),
    .B(_03850_),
    .X(_03851_));
 sky130_fd_sc_hd__a21boi_1 _20624_ (.A1(_03844_),
    .A2(_03846_),
    .B1_N(_03845_),
    .Y(_03852_));
 sky130_fd_sc_hd__xnor2_1 _20625_ (.A(_03851_),
    .B(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hd__a22o_1 _20626_ (.A1(\rbzero.texV[-3] ),
    .A2(_03814_),
    .B1(_03819_),
    .B2(_03853_),
    .X(_01608_));
 sky130_fd_sc_hd__or2_1 _20627_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .X(_03854_));
 sky130_fd_sc_hd__nand2_1 _20628_ (.A(\rbzero.traced_texa[-2] ),
    .B(\rbzero.texV[-2] ),
    .Y(_03855_));
 sky130_fd_sc_hd__o21ai_1 _20629_ (.A1(_03849_),
    .A2(_03852_),
    .B1(_03850_),
    .Y(_03856_));
 sky130_fd_sc_hd__nand3_1 _20630_ (.A(_03854_),
    .B(_03855_),
    .C(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__a21o_1 _20631_ (.A1(_03854_),
    .A2(_03855_),
    .B1(_03856_),
    .X(_03858_));
 sky130_fd_sc_hd__a32o_1 _20632_ (.A1(_03734_),
    .A2(_03857_),
    .A3(_03858_),
    .B1(_03740_),
    .B2(\rbzero.texV[-2] ),
    .X(_01609_));
 sky130_fd_sc_hd__nor2_1 _20633_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .Y(_03859_));
 sky130_fd_sc_hd__and2_1 _20634_ (.A(\rbzero.traced_texa[-1] ),
    .B(\rbzero.texV[-1] ),
    .X(_03860_));
 sky130_fd_sc_hd__or2_1 _20635_ (.A(_03859_),
    .B(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__a21boi_1 _20636_ (.A1(_03854_),
    .A2(_03856_),
    .B1_N(_03855_),
    .Y(_03862_));
 sky130_fd_sc_hd__xor2_1 _20637_ (.A(_03861_),
    .B(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__a22o_1 _20638_ (.A1(\rbzero.texV[-1] ),
    .A2(_03814_),
    .B1(_03819_),
    .B2(_03863_),
    .X(_01610_));
 sky130_fd_sc_hd__nor2_1 _20639_ (.A(_03861_),
    .B(_03862_),
    .Y(_03864_));
 sky130_fd_sc_hd__or2_1 _20640_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .X(_03865_));
 sky130_fd_sc_hd__nand2_1 _20641_ (.A(\rbzero.traced_texa[0] ),
    .B(\rbzero.texV[0] ),
    .Y(_03866_));
 sky130_fd_sc_hd__o211a_1 _20642_ (.A1(_03860_),
    .A2(_03864_),
    .B1(_03865_),
    .C1(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__inv_2 _20643_ (.A(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__a211o_1 _20644_ (.A1(_03865_),
    .A2(_03866_),
    .B1(_03860_),
    .C1(_03864_),
    .X(_03869_));
 sky130_fd_sc_hd__a32o_1 _20645_ (.A1(_03734_),
    .A2(_03868_),
    .A3(_03869_),
    .B1(_03740_),
    .B2(\rbzero.texV[0] ),
    .X(_01611_));
 sky130_fd_sc_hd__or2_1 _20646_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .X(_03870_));
 sky130_fd_sc_hd__nand2_1 _20647_ (.A(\rbzero.traced_texa[1] ),
    .B(\rbzero.texV[1] ),
    .Y(_03871_));
 sky130_fd_sc_hd__nand2_1 _20648_ (.A(_03866_),
    .B(_03868_),
    .Y(_03872_));
 sky130_fd_sc_hd__a21o_1 _20649_ (.A1(_03870_),
    .A2(_03871_),
    .B1(_03872_),
    .X(_03873_));
 sky130_fd_sc_hd__and3_1 _20650_ (.A(_03870_),
    .B(_03871_),
    .C(_03872_),
    .X(_03874_));
 sky130_fd_sc_hd__inv_2 _20651_ (.A(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__a32o_1 _20652_ (.A1(_03734_),
    .A2(_03873_),
    .A3(_03875_),
    .B1(_03740_),
    .B2(\rbzero.texV[1] ),
    .X(_01612_));
 sky130_fd_sc_hd__or2_1 _20653_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .X(_03876_));
 sky130_fd_sc_hd__nand2_1 _20654_ (.A(\rbzero.traced_texa[2] ),
    .B(\rbzero.texV[2] ),
    .Y(_03877_));
 sky130_fd_sc_hd__nand2_1 _20655_ (.A(_03871_),
    .B(_03875_),
    .Y(_03878_));
 sky130_fd_sc_hd__a21o_1 _20656_ (.A1(_03876_),
    .A2(_03877_),
    .B1(_03878_),
    .X(_03879_));
 sky130_fd_sc_hd__and3_1 _20657_ (.A(_03876_),
    .B(_03877_),
    .C(_03878_),
    .X(_03880_));
 sky130_fd_sc_hd__inv_2 _20658_ (.A(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__a32o_1 _20659_ (.A1(_03734_),
    .A2(_03879_),
    .A3(_03881_),
    .B1(_03740_),
    .B2(\rbzero.texV[2] ),
    .X(_01613_));
 sky130_fd_sc_hd__or2_1 _20660_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .X(_03882_));
 sky130_fd_sc_hd__nand2_1 _20661_ (.A(\rbzero.traced_texa[3] ),
    .B(\rbzero.texV[3] ),
    .Y(_03883_));
 sky130_fd_sc_hd__nand2_1 _20662_ (.A(_03877_),
    .B(_03881_),
    .Y(_03884_));
 sky130_fd_sc_hd__and3_1 _20663_ (.A(_03882_),
    .B(_03883_),
    .C(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__inv_2 _20664_ (.A(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__a21o_1 _20665_ (.A1(_03882_),
    .A2(_03883_),
    .B1(_03884_),
    .X(_03887_));
 sky130_fd_sc_hd__a32o_1 _20666_ (.A1(_03734_),
    .A2(_03886_),
    .A3(_03887_),
    .B1(_03740_),
    .B2(\rbzero.texV[3] ),
    .X(_01614_));
 sky130_fd_sc_hd__or2_1 _20667_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .X(_03888_));
 sky130_fd_sc_hd__nand2_1 _20668_ (.A(\rbzero.traced_texa[4] ),
    .B(\rbzero.texV[4] ),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2_1 _20669_ (.A(_03883_),
    .B(_03886_),
    .Y(_03890_));
 sky130_fd_sc_hd__a21o_1 _20670_ (.A1(_03888_),
    .A2(_03889_),
    .B1(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__nand3_1 _20671_ (.A(_03888_),
    .B(_03889_),
    .C(_03890_),
    .Y(_03892_));
 sky130_fd_sc_hd__a32o_1 _20672_ (.A1(_09732_),
    .A2(_03891_),
    .A3(_03892_),
    .B1(_03740_),
    .B2(\rbzero.texV[4] ),
    .X(_01615_));
 sky130_fd_sc_hd__a21boi_1 _20673_ (.A1(_03888_),
    .A2(_03890_),
    .B1_N(_03889_),
    .Y(_03893_));
 sky130_fd_sc_hd__nor2_1 _20674_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_03894_));
 sky130_fd_sc_hd__nand2_1 _20675_ (.A(\rbzero.traced_texa[5] ),
    .B(\rbzero.texV[5] ),
    .Y(_03895_));
 sky130_fd_sc_hd__and2b_1 _20676_ (.A_N(_03894_),
    .B(_03895_),
    .X(_03896_));
 sky130_fd_sc_hd__xnor2_1 _20677_ (.A(_03893_),
    .B(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__a22o_1 _20678_ (.A1(\rbzero.texV[5] ),
    .A2(_03814_),
    .B1(_03819_),
    .B2(_03897_),
    .X(_01616_));
 sky130_fd_sc_hd__or2_1 _20679_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .X(_03898_));
 sky130_fd_sc_hd__nand2_1 _20680_ (.A(\rbzero.traced_texa[6] ),
    .B(\rbzero.texV[6] ),
    .Y(_03899_));
 sky130_fd_sc_hd__nand2_1 _20681_ (.A(_03898_),
    .B(_03899_),
    .Y(_03900_));
 sky130_fd_sc_hd__o21ai_1 _20682_ (.A1(_03893_),
    .A2(_03894_),
    .B1(_03895_),
    .Y(_03901_));
 sky130_fd_sc_hd__xnor2_1 _20683_ (.A(_03900_),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__a22o_1 _20684_ (.A1(\rbzero.texV[6] ),
    .A2(_03814_),
    .B1(_03819_),
    .B2(_03902_),
    .X(_01617_));
 sky130_fd_sc_hd__nor2_1 _20685_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_03903_));
 sky130_fd_sc_hd__nand2_1 _20686_ (.A(\rbzero.traced_texa[7] ),
    .B(\rbzero.texV[7] ),
    .Y(_03904_));
 sky130_fd_sc_hd__and2b_1 _20687_ (.A_N(_03903_),
    .B(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__a21boi_1 _20688_ (.A1(_03898_),
    .A2(_03901_),
    .B1_N(_03899_),
    .Y(_03906_));
 sky130_fd_sc_hd__xnor2_1 _20689_ (.A(_03905_),
    .B(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__a22o_1 _20690_ (.A1(\rbzero.texV[7] ),
    .A2(_03814_),
    .B1(_03819_),
    .B2(_03907_),
    .X(_01618_));
 sky130_fd_sc_hd__or2_1 _20691_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .X(_03908_));
 sky130_fd_sc_hd__nand2_1 _20692_ (.A(\rbzero.traced_texa[8] ),
    .B(\rbzero.texV[8] ),
    .Y(_03909_));
 sky130_fd_sc_hd__o21ai_1 _20693_ (.A1(_03903_),
    .A2(_03906_),
    .B1(_03904_),
    .Y(_03910_));
 sky130_fd_sc_hd__a21o_1 _20694_ (.A1(_03908_),
    .A2(_03909_),
    .B1(_03910_),
    .X(_03911_));
 sky130_fd_sc_hd__nand3_1 _20695_ (.A(_03908_),
    .B(_03909_),
    .C(_03910_),
    .Y(_03912_));
 sky130_fd_sc_hd__a32o_1 _20696_ (.A1(_09732_),
    .A2(_03911_),
    .A3(_03912_),
    .B1(_03740_),
    .B2(\rbzero.texV[8] ),
    .X(_01619_));
 sky130_fd_sc_hd__or2_1 _20697_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .X(_03913_));
 sky130_fd_sc_hd__nand2_1 _20698_ (.A(\rbzero.traced_texa[9] ),
    .B(\rbzero.texV[9] ),
    .Y(_03914_));
 sky130_fd_sc_hd__a21o_1 _20699_ (.A1(\rbzero.traced_texa[8] ),
    .A2(\rbzero.texV[8] ),
    .B1(_03910_),
    .X(_03915_));
 sky130_fd_sc_hd__a22o_1 _20700_ (.A1(_03913_),
    .A2(_03914_),
    .B1(_03915_),
    .B2(_03908_),
    .X(_03916_));
 sky130_fd_sc_hd__nand4_1 _20701_ (.A(_03908_),
    .B(_03913_),
    .C(_03914_),
    .D(_03915_),
    .Y(_03917_));
 sky130_fd_sc_hd__a32o_1 _20702_ (.A1(_09732_),
    .A2(_03916_),
    .A3(_03917_),
    .B1(_03740_),
    .B2(\rbzero.texV[9] ),
    .X(_01620_));
 sky130_fd_sc_hd__xnor2_1 _20703_ (.A(\rbzero.traced_texa[10] ),
    .B(\rbzero.texV[10] ),
    .Y(_03918_));
 sky130_fd_sc_hd__and3_1 _20704_ (.A(_03914_),
    .B(_03917_),
    .C(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__a21oi_1 _20705_ (.A1(_03914_),
    .A2(_03917_),
    .B1(_03918_),
    .Y(_03920_));
 sky130_fd_sc_hd__nor2_1 _20706_ (.A(_03919_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__a22o_1 _20707_ (.A1(\rbzero.texV[10] ),
    .A2(_03814_),
    .B1(_03819_),
    .B2(_03921_),
    .X(_01621_));
 sky130_fd_sc_hd__o21ai_1 _20708_ (.A1(_04436_),
    .A2(_08141_),
    .B1(_04437_),
    .Y(_03922_));
 sky130_fd_sc_hd__nand2_1 _20709_ (.A(_04437_),
    .B(_09729_),
    .Y(_03923_));
 sky130_fd_sc_hd__a21o_1 _20710_ (.A1(_05050_),
    .A2(_03923_),
    .B1(_08045_),
    .X(_03924_));
 sky130_fd_sc_hd__mux2_1 _20711_ (.A0(_03922_),
    .A1(_04437_),
    .S(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__and2_1 _20712_ (.A(_04442_),
    .B(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__clkbuf_1 _20713_ (.A(_03926_),
    .X(_01622_));
 sky130_fd_sc_hd__nand2_1 _20714_ (.A(_04436_),
    .B(_04437_),
    .Y(_03927_));
 sky130_fd_sc_hd__o211a_1 _20715_ (.A1(_03927_),
    .A2(_03924_),
    .B1(_04442_),
    .C1(_04430_),
    .X(_01623_));
 sky130_fd_sc_hd__nor2_1 _20716_ (.A(_03927_),
    .B(_03924_),
    .Y(_03928_));
 sky130_fd_sc_hd__a21oi_1 _20717_ (.A1(_04429_),
    .A2(_03928_),
    .B1(_08136_),
    .Y(_03929_));
 sky130_fd_sc_hd__o21a_1 _20718_ (.A1(_04429_),
    .A2(_03928_),
    .B1(_03929_),
    .X(_01624_));
 sky130_fd_sc_hd__a21boi_1 _20719_ (.A1(_04429_),
    .A2(_04436_),
    .B1_N(\rbzero.trace_state[3] ),
    .Y(_03930_));
 sky130_fd_sc_hd__o31a_1 _20720_ (.A1(_08405_),
    .A2(_03924_),
    .A3(_03930_),
    .B1(_01633_),
    .X(_01625_));
 sky130_fd_sc_hd__and2_2 _20721_ (.A(_08117_),
    .B(clknet_1_0__leaf__05700_),
    .X(_03931_));
 sky130_fd_sc_hd__buf_1 _20722_ (.A(_03931_),
    .X(_01626_));
 sky130_fd_sc_hd__and2_2 _20723_ (.A(_03728_),
    .B(clknet_1_0__leaf__05761_),
    .X(_03932_));
 sky130_fd_sc_hd__buf_1 _20724_ (.A(_03932_),
    .X(_01627_));
 sky130_fd_sc_hd__and2_2 _20725_ (.A(_03728_),
    .B(clknet_1_0__leaf__05820_),
    .X(_03933_));
 sky130_fd_sc_hd__buf_1 _20726_ (.A(_03933_),
    .X(_01628_));
 sky130_fd_sc_hd__and2_2 _20727_ (.A(_03728_),
    .B(clknet_1_1__leaf__05879_),
    .X(_03934_));
 sky130_fd_sc_hd__buf_1 _20728_ (.A(_03934_),
    .X(_01629_));
 sky130_fd_sc_hd__and2_2 _20729_ (.A(_03728_),
    .B(clknet_1_0__leaf__05938_),
    .X(_03935_));
 sky130_fd_sc_hd__buf_1 _20730_ (.A(_03935_),
    .X(_01630_));
 sky130_fd_sc_hd__and2_2 _20731_ (.A(_03728_),
    .B(clknet_1_1__leaf__05993_),
    .X(_03936_));
 sky130_fd_sc_hd__buf_1 _20732_ (.A(_03936_),
    .X(_01631_));
 sky130_fd_sc_hd__nor2_1 _20733_ (.A(\rbzero.hsync ),
    .B(net63),
    .Y(_01632_));
 sky130_fd_sc_hd__buf_2 _20734_ (.A(_09749_),
    .X(_03937_));
 sky130_fd_sc_hd__a22o_1 _20735_ (.A1(\rbzero.traced_texVinit[0] ),
    .A2(_09759_),
    .B1(_03937_),
    .B2(_09111_),
    .X(_01634_));
 sky130_fd_sc_hd__a22o_1 _20736_ (.A1(\rbzero.traced_texVinit[1] ),
    .A2(_09759_),
    .B1(_03937_),
    .B2(_09105_),
    .X(_01635_));
 sky130_fd_sc_hd__a22o_1 _20737_ (.A1(\rbzero.traced_texVinit[2] ),
    .A2(_09759_),
    .B1(_03937_),
    .B2(_09101_),
    .X(_01636_));
 sky130_fd_sc_hd__a22o_1 _20738_ (.A1(\rbzero.traced_texVinit[3] ),
    .A2(_09759_),
    .B1(_03937_),
    .B2(_09227_),
    .X(_01637_));
 sky130_fd_sc_hd__a22o_1 _20739_ (.A1(\rbzero.traced_texVinit[4] ),
    .A2(_09759_),
    .B1(_03937_),
    .B2(_09347_),
    .X(_01638_));
 sky130_fd_sc_hd__a22o_1 _20740_ (.A1(\rbzero.traced_texVinit[5] ),
    .A2(_09759_),
    .B1(_03937_),
    .B2(_09868_),
    .X(_01639_));
 sky130_fd_sc_hd__a22o_1 _20741_ (.A1(\rbzero.traced_texVinit[6] ),
    .A2(_09759_),
    .B1(_03937_),
    .B2(_09593_),
    .X(_01640_));
 sky130_fd_sc_hd__a22o_1 _20742_ (.A1(\rbzero.traced_texVinit[7] ),
    .A2(_09759_),
    .B1(_03937_),
    .B2(_09721_),
    .X(_01641_));
 sky130_fd_sc_hd__a22o_1 _20743_ (.A1(\rbzero.traced_texVinit[8] ),
    .A2(_09759_),
    .B1(_03937_),
    .B2(_10010_),
    .X(_01642_));
 sky130_fd_sc_hd__a22o_1 _20744_ (.A1(\rbzero.traced_texVinit[9] ),
    .A2(_02606_),
    .B1(_03937_),
    .B2(_10126_),
    .X(_01643_));
 sky130_fd_sc_hd__a22o_1 _20745_ (.A1(\rbzero.traced_texVinit[10] ),
    .A2(_02606_),
    .B1(_02557_),
    .B2(_10258_),
    .X(_01644_));
 sky130_fd_sc_hd__nor2_1 _20746_ (.A(\gpout0.clk_div[0] ),
    .B(net63),
    .Y(_01645_));
 sky130_fd_sc_hd__nand2_1 _20747_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .Y(_03938_));
 sky130_fd_sc_hd__or2_1 _20748_ (.A(\gpout0.clk_div[0] ),
    .B(\gpout0.clk_div[1] ),
    .X(_03939_));
 sky130_fd_sc_hd__and3_1 _20749_ (.A(_03728_),
    .B(_03938_),
    .C(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__clkbuf_1 _20750_ (.A(_03940_),
    .X(_01646_));
 sky130_fd_sc_hd__or2_1 _20751_ (.A(\rbzero.debug_overlay.vplaneX[-9] ),
    .B(\rbzero.wall_tracer.rayAddendX[-9] ),
    .X(_03941_));
 sky130_fd_sc_hd__and3_1 _20752_ (.A(_09749_),
    .B(_02514_),
    .C(_03941_),
    .X(_03942_));
 sky130_fd_sc_hd__a21o_1 _20753_ (.A1(\rbzero.wall_tracer.rayAddendX[-9] ),
    .A2(_09746_),
    .B1(_03942_),
    .X(_01647_));
 sky130_fd_sc_hd__nor2_1 _20754_ (.A(_02516_),
    .B(_02515_),
    .Y(_03943_));
 sky130_fd_sc_hd__xnor2_1 _20755_ (.A(_02514_),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__a22o_1 _20756_ (.A1(\rbzero.wall_tracer.rayAddendX[-8] ),
    .A2(_02606_),
    .B1(_02557_),
    .B2(_03944_),
    .X(_01648_));
 sky130_fd_sc_hd__and2b_1 _20757_ (.A_N(_02513_),
    .B(_02518_),
    .X(_03945_));
 sky130_fd_sc_hd__xnor2_1 _20758_ (.A(_02517_),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__a22o_1 _20759_ (.A1(\rbzero.wall_tracer.rayAddendX[-7] ),
    .A2(_02606_),
    .B1(_02557_),
    .B2(_03946_),
    .X(_01649_));
 sky130_fd_sc_hd__xnor2_1 _20760_ (.A(_05120_),
    .B(\rbzero.wall_tracer.rayAddendX[-6] ),
    .Y(_03947_));
 sky130_fd_sc_hd__xnor2_1 _20761_ (.A(_02519_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__a22o_1 _20762_ (.A1(\rbzero.wall_tracer.rayAddendX[-6] ),
    .A2(_02606_),
    .B1(_02557_),
    .B2(_03948_),
    .X(_01650_));
 sky130_fd_sc_hd__or2_1 _20763_ (.A(\rbzero.debug_overlay.vplaneY[-9] ),
    .B(\rbzero.wall_tracer.rayAddendY[-9] ),
    .X(_03949_));
 sky130_fd_sc_hd__and3_1 _20764_ (.A(_09749_),
    .B(_02747_),
    .C(_03949_),
    .X(_03950_));
 sky130_fd_sc_hd__a21o_1 _20765_ (.A1(\rbzero.wall_tracer.rayAddendY[-9] ),
    .A2(_09746_),
    .B1(_03950_),
    .X(_01651_));
 sky130_fd_sc_hd__nor2_1 _20766_ (.A(_02749_),
    .B(_02748_),
    .Y(_03951_));
 sky130_fd_sc_hd__xnor2_1 _20767_ (.A(_02747_),
    .B(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__a22o_1 _20768_ (.A1(\rbzero.wall_tracer.rayAddendY[-8] ),
    .A2(_02606_),
    .B1(_02557_),
    .B2(_03952_),
    .X(_01652_));
 sky130_fd_sc_hd__and2b_1 _20769_ (.A_N(_02746_),
    .B(_02751_),
    .X(_03953_));
 sky130_fd_sc_hd__xnor2_1 _20770_ (.A(_02750_),
    .B(_03953_),
    .Y(_03954_));
 sky130_fd_sc_hd__a22o_1 _20771_ (.A1(\rbzero.wall_tracer.rayAddendY[-7] ),
    .A2(_02606_),
    .B1(_02557_),
    .B2(_03954_),
    .X(_01653_));
 sky130_fd_sc_hd__xnor2_1 _20772_ (.A(_05129_),
    .B(\rbzero.wall_tracer.rayAddendY[-6] ),
    .Y(_03955_));
 sky130_fd_sc_hd__xnor2_1 _20773_ (.A(_02752_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__a22o_1 _20774_ (.A1(\rbzero.wall_tracer.rayAddendY[-6] ),
    .A2(_02606_),
    .B1(_02557_),
    .B2(_03956_),
    .X(_01654_));
 sky130_fd_sc_hd__nor2_1 _20775_ (.A(\gpout1.clk_div[0] ),
    .B(net63),
    .Y(_01655_));
 sky130_fd_sc_hd__nand2_1 _20776_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .Y(_03957_));
 sky130_fd_sc_hd__or2_1 _20777_ (.A(\gpout1.clk_div[0] ),
    .B(\gpout1.clk_div[1] ),
    .X(_03958_));
 sky130_fd_sc_hd__and3_1 _20778_ (.A(_03728_),
    .B(_03957_),
    .C(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__clkbuf_1 _20779_ (.A(_03959_),
    .X(_01656_));
 sky130_fd_sc_hd__nor2_1 _20780_ (.A(\gpout2.clk_div[0] ),
    .B(net63),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_1 _20781_ (.A(\gpout2.clk_div[1] ),
    .B(\gpout2.clk_div[0] ),
    .Y(_03960_));
 sky130_fd_sc_hd__or2_1 _20782_ (.A(\gpout2.clk_div[1] ),
    .B(\gpout2.clk_div[0] ),
    .X(_03961_));
 sky130_fd_sc_hd__and3_1 _20783_ (.A(_03110_),
    .B(_03960_),
    .C(_03961_),
    .X(_03962_));
 sky130_fd_sc_hd__clkbuf_1 _20784_ (.A(_03962_),
    .X(_01658_));
 sky130_fd_sc_hd__nor2_1 _20785_ (.A(\gpout3.clk_div[0] ),
    .B(net63),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_1 _20786_ (.A(\gpout3.clk_div[0] ),
    .B(\gpout3.clk_div[1] ),
    .Y(_03963_));
 sky130_fd_sc_hd__or2_1 _20787_ (.A(\gpout3.clk_div[0] ),
    .B(\gpout3.clk_div[1] ),
    .X(_03964_));
 sky130_fd_sc_hd__and3_1 _20788_ (.A(_03110_),
    .B(_03963_),
    .C(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__clkbuf_1 _20789_ (.A(_03965_),
    .X(_01660_));
 sky130_fd_sc_hd__nor2_1 _20790_ (.A(\gpout4.clk_div[0] ),
    .B(net63),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_1 _20791_ (.A(\gpout4.clk_div[0] ),
    .B(\gpout4.clk_div[1] ),
    .Y(_03966_));
 sky130_fd_sc_hd__or2_1 _20792_ (.A(\gpout4.clk_div[0] ),
    .B(\gpout4.clk_div[1] ),
    .X(_03967_));
 sky130_fd_sc_hd__and3_1 _20793_ (.A(_03110_),
    .B(_03966_),
    .C(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__clkbuf_1 _20794_ (.A(_03968_),
    .X(_01662_));
 sky130_fd_sc_hd__dfxtp_4 _20795_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00000_),
    .Q(\rbzero.wall_tracer.rcp_sel[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20796_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00001_),
    .Q(\rbzero.wall_tracer.rcp_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20797_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00386_),
    .Q(\rbzero.wall_tracer.mapY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20798_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00387_),
    .Q(\rbzero.wall_tracer.mapY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20799_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00388_),
    .Q(\rbzero.wall_tracer.mapY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20800_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00389_),
    .Q(\rbzero.wall_tracer.mapY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20801_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00390_),
    .Q(\rbzero.wall_tracer.mapY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20802_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00391_),
    .Q(\rbzero.wall_tracer.stepDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20803_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00392_),
    .Q(\rbzero.wall_tracer.stepDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20804_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00393_),
    .Q(\rbzero.wall_tracer.stepDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20805_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00394_),
    .Q(\rbzero.wall_tracer.stepDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20806_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00395_),
    .Q(\rbzero.wall_tracer.stepDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20807_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00396_),
    .Q(\rbzero.wall_tracer.stepDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20808_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00397_),
    .Q(\rbzero.wall_tracer.stepDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20809_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00398_),
    .Q(\rbzero.wall_tracer.stepDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20810_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00399_),
    .Q(\rbzero.wall_tracer.stepDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20811_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00400_),
    .Q(\rbzero.wall_tracer.stepDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20812_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00401_),
    .Q(\rbzero.wall_tracer.stepDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20813_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00402_),
    .Q(\rbzero.wall_tracer.stepDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20814_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00403_),
    .Q(\rbzero.wall_tracer.stepDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20815_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00404_),
    .Q(\rbzero.wall_tracer.stepDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20816_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00405_),
    .Q(\rbzero.wall_tracer.stepDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20817_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00406_),
    .Q(\rbzero.wall_tracer.stepDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20818_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00407_),
    .Q(\rbzero.wall_tracer.stepDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20819_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00408_),
    .Q(\rbzero.wall_tracer.stepDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20820_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00409_),
    .Q(\rbzero.wall_tracer.stepDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20821_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00410_),
    .Q(\rbzero.wall_tracer.stepDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20822_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00411_),
    .Q(\rbzero.wall_tracer.stepDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20823_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00412_),
    .Q(\rbzero.wall_tracer.stepDistY[10] ));
 sky130_fd_sc_hd__dfxtp_4 _20824_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00413_),
    .Q(\rbzero.wall_tracer.visualWallDist[-11] ));
 sky130_fd_sc_hd__dfxtp_4 _20825_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00414_),
    .Q(\rbzero.wall_tracer.visualWallDist[-10] ));
 sky130_fd_sc_hd__dfxtp_2 _20826_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00415_),
    .Q(\rbzero.wall_tracer.visualWallDist[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20827_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00416_),
    .Q(\rbzero.wall_tracer.visualWallDist[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20828_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00417_),
    .Q(\rbzero.wall_tracer.visualWallDist[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20829_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00418_),
    .Q(\rbzero.wall_tracer.visualWallDist[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20830_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00419_),
    .Q(\rbzero.wall_tracer.visualWallDist[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20831_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00420_),
    .Q(\rbzero.wall_tracer.visualWallDist[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20832_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00421_),
    .Q(\rbzero.wall_tracer.visualWallDist[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _20833_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00422_),
    .Q(\rbzero.wall_tracer.visualWallDist[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _20834_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00423_),
    .Q(\rbzero.wall_tracer.visualWallDist[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _20835_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00424_),
    .Q(\rbzero.wall_tracer.visualWallDist[0] ));
 sky130_fd_sc_hd__dfxtp_4 _20836_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00425_),
    .Q(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__dfxtp_4 _20837_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00426_),
    .Q(\rbzero.wall_tracer.visualWallDist[2] ));
 sky130_fd_sc_hd__dfxtp_4 _20838_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00427_),
    .Q(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__dfxtp_4 _20839_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00428_),
    .Q(\rbzero.wall_tracer.visualWallDist[4] ));
 sky130_fd_sc_hd__dfxtp_4 _20840_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00429_),
    .Q(\rbzero.wall_tracer.visualWallDist[5] ));
 sky130_fd_sc_hd__dfxtp_4 _20841_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00430_),
    .Q(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__dfxtp_4 _20842_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00431_),
    .Q(\rbzero.wall_tracer.visualWallDist[7] ));
 sky130_fd_sc_hd__dfxtp_4 _20843_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00432_),
    .Q(\rbzero.wall_tracer.visualWallDist[8] ));
 sky130_fd_sc_hd__dfxtp_4 _20844_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00433_),
    .Q(\rbzero.wall_tracer.visualWallDist[9] ));
 sky130_fd_sc_hd__dfxtp_4 _20845_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00434_),
    .Q(\rbzero.wall_tracer.visualWallDist[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20846_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00435_),
    .Q(\rbzero.wall_tracer.stepDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20847_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00436_),
    .Q(\rbzero.wall_tracer.stepDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20848_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00437_),
    .Q(\rbzero.wall_tracer.stepDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20849_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00438_),
    .Q(\rbzero.wall_tracer.stepDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20850_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00439_),
    .Q(\rbzero.wall_tracer.stepDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20851_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00440_),
    .Q(\rbzero.wall_tracer.stepDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20852_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00441_),
    .Q(\rbzero.wall_tracer.stepDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_2 _20853_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00442_),
    .Q(\rbzero.wall_tracer.stepDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _20854_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00443_),
    .Q(\rbzero.wall_tracer.stepDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20855_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00444_),
    .Q(\rbzero.wall_tracer.stepDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20856_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00445_),
    .Q(\rbzero.wall_tracer.stepDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20857_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00446_),
    .Q(\rbzero.wall_tracer.stepDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20858_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00447_),
    .Q(\rbzero.wall_tracer.stepDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20859_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00448_),
    .Q(\rbzero.wall_tracer.stepDistX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20860_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00449_),
    .Q(\rbzero.wall_tracer.stepDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20861_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00450_),
    .Q(\rbzero.wall_tracer.stepDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20862_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00451_),
    .Q(\rbzero.wall_tracer.stepDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20863_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00452_),
    .Q(\rbzero.wall_tracer.stepDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20864_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00453_),
    .Q(\rbzero.wall_tracer.stepDistX[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20865_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00454_),
    .Q(\rbzero.wall_tracer.stepDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20866_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00455_),
    .Q(\rbzero.wall_tracer.stepDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20867_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00456_),
    .Q(\rbzero.wall_tracer.stepDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20868_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00457_),
    .Q(\reg_rgb[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20869_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00458_),
    .Q(\reg_rgb[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20870_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00459_),
    .Q(\reg_rgb[14] ));
 sky130_fd_sc_hd__dfxtp_1 _20871_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00460_),
    .Q(\reg_rgb[15] ));
 sky130_fd_sc_hd__dfxtp_1 _20872_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00461_),
    .Q(\reg_rgb[22] ));
 sky130_fd_sc_hd__dfxtp_1 _20873_ (.CLK(clknet_leaf_43_i_clk),
    .D(_00462_),
    .Q(\reg_rgb[23] ));
 sky130_fd_sc_hd__dfxtp_4 _20874_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00463_),
    .Q(\rbzero.wall_hot[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20875_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00464_),
    .Q(\rbzero.wall_hot[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20876_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00465_),
    .Q(\rbzero.side_hot ));
 sky130_fd_sc_hd__dfxtp_1 _20877_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00466_),
    .Q(\rbzero.texu_hot[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20878_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00467_),
    .Q(\rbzero.texu_hot[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20879_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00468_),
    .Q(\rbzero.texu_hot[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20880_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00469_),
    .Q(\rbzero.texu_hot[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20881_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00470_),
    .Q(\rbzero.texu_hot[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20882_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00471_),
    .Q(\rbzero.texu_hot[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20883_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00472_),
    .Q(\gpout0.hpos[0] ));
 sky130_fd_sc_hd__dfxtp_4 _20884_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00473_),
    .Q(\gpout0.hpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20885_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00474_),
    .Q(\gpout0.hpos[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20886_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00475_),
    .Q(\gpout0.hpos[3] ));
 sky130_fd_sc_hd__dfxtp_4 _20887_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00476_),
    .Q(\gpout0.hpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20888_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00477_),
    .Q(\gpout0.hpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20889_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00478_),
    .Q(\gpout0.hpos[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20890_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00479_),
    .Q(\gpout0.hpos[7] ));
 sky130_fd_sc_hd__dfxtp_4 _20891_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00480_),
    .Q(\gpout0.hpos[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20892_ (.CLK(clknet_leaf_44_i_clk),
    .D(_00481_),
    .Q(\gpout0.hpos[9] ));
 sky130_fd_sc_hd__dfxtp_4 _20893_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00482_),
    .Q(\rbzero.row_render.side ));
 sky130_fd_sc_hd__dfxtp_1 _20894_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00483_),
    .Q(\rbzero.row_render.size[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20895_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00484_),
    .Q(\rbzero.row_render.size[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20896_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00485_),
    .Q(\rbzero.row_render.size[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20897_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00486_),
    .Q(\rbzero.row_render.size[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20898_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00487_),
    .Q(\rbzero.row_render.size[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20899_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00488_),
    .Q(\rbzero.row_render.size[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20900_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00489_),
    .Q(\rbzero.row_render.size[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20901_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00490_),
    .Q(\rbzero.row_render.size[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20902_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00491_),
    .Q(\rbzero.row_render.size[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20903_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00492_),
    .Q(\rbzero.row_render.size[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20904_ (.CLK(clknet_leaf_41_i_clk),
    .D(_00493_),
    .Q(\rbzero.row_render.size[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20905_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00494_),
    .Q(\rbzero.row_render.texu[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20906_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00495_),
    .Q(\rbzero.row_render.texu[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20907_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00496_),
    .Q(\rbzero.row_render.texu[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20908_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00497_),
    .Q(\rbzero.row_render.texu[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20909_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00498_),
    .Q(\rbzero.row_render.texu[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20910_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00499_),
    .Q(\rbzero.traced_texa[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20911_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00500_),
    .Q(\rbzero.traced_texa[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20912_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00501_),
    .Q(\rbzero.traced_texa[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20913_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00502_),
    .Q(\rbzero.traced_texa[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20914_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00503_),
    .Q(\rbzero.traced_texa[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20915_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00504_),
    .Q(\rbzero.traced_texa[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20916_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00505_),
    .Q(\rbzero.traced_texa[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20917_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00506_),
    .Q(\rbzero.traced_texa[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20918_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00507_),
    .Q(\rbzero.traced_texa[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20919_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00508_),
    .Q(\rbzero.traced_texa[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20920_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00509_),
    .Q(\rbzero.traced_texa[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20921_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00510_),
    .Q(\rbzero.traced_texa[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20922_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00511_),
    .Q(\rbzero.traced_texa[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20923_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00512_),
    .Q(\rbzero.traced_texa[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20924_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00513_),
    .Q(\rbzero.traced_texa[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20925_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00514_),
    .Q(\rbzero.traced_texa[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20926_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00515_),
    .Q(\rbzero.traced_texa[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20927_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00516_),
    .Q(\rbzero.traced_texa[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20928_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00517_),
    .Q(\rbzero.traced_texa[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20929_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00518_),
    .Q(\rbzero.traced_texa[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20930_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00519_),
    .Q(\rbzero.traced_texa[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20931_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00520_),
    .Q(\rbzero.traced_texa[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20932_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00521_),
    .Q(\rbzero.row_render.wall[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20933_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00522_),
    .Q(\rbzero.row_render.wall[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20934_ (.CLK(clknet_leaf_45_i_clk),
    .D(_00523_),
    .Q(\rbzero.wall_tracer.mapX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20935_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00524_),
    .Q(\rbzero.wall_tracer.mapX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20936_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00525_),
    .Q(\rbzero.wall_tracer.mapX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20937_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00526_),
    .Q(\rbzero.wall_tracer.mapX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20938_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00527_),
    .Q(\rbzero.wall_tracer.mapX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20939_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00528_),
    .Q(\rbzero.wall_tracer.trackDistX[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20940_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00529_),
    .Q(\rbzero.wall_tracer.trackDistX[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20941_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00530_),
    .Q(\rbzero.wall_tracer.trackDistX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20942_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00531_),
    .Q(\rbzero.wall_tracer.trackDistX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20943_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00532_),
    .Q(\rbzero.wall_tracer.trackDistX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20944_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00533_),
    .Q(\rbzero.wall_tracer.trackDistX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20945_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00534_),
    .Q(\rbzero.wall_tracer.trackDistX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20946_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00535_),
    .Q(\rbzero.wall_tracer.trackDistX[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20947_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00536_),
    .Q(\rbzero.wall_tracer.trackDistX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20948_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00537_),
    .Q(\rbzero.wall_tracer.trackDistX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20949_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00538_),
    .Q(\rbzero.wall_tracer.trackDistX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20950_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00539_),
    .Q(\rbzero.wall_tracer.trackDistX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20951_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00540_),
    .Q(\rbzero.wall_tracer.trackDistX[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20952_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00541_),
    .Q(\rbzero.wall_tracer.trackDistX[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20953_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00542_),
    .Q(\rbzero.wall_tracer.trackDistX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20954_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00543_),
    .Q(\rbzero.wall_tracer.trackDistX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20955_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00544_),
    .Q(\rbzero.wall_tracer.trackDistX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20956_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00545_),
    .Q(\rbzero.wall_tracer.trackDistX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20957_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00546_),
    .Q(\rbzero.wall_tracer.trackDistX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20958_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00547_),
    .Q(\rbzero.wall_tracer.trackDistX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20959_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00548_),
    .Q(\rbzero.wall_tracer.trackDistX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20960_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00549_),
    .Q(\rbzero.wall_tracer.trackDistX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20961_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00550_),
    .Q(\rbzero.wall_tracer.trackDistY[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _20962_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00551_),
    .Q(\rbzero.wall_tracer.trackDistY[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _20963_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00552_),
    .Q(\rbzero.wall_tracer.trackDistY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _20964_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00553_),
    .Q(\rbzero.wall_tracer.trackDistY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _20965_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00554_),
    .Q(\rbzero.wall_tracer.trackDistY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _20966_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00555_),
    .Q(\rbzero.wall_tracer.trackDistY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _20967_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00556_),
    .Q(\rbzero.wall_tracer.trackDistY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _20968_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00557_),
    .Q(\rbzero.wall_tracer.trackDistY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _20969_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00558_),
    .Q(\rbzero.wall_tracer.trackDistY[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _20970_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00559_),
    .Q(\rbzero.wall_tracer.trackDistY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _20971_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00560_),
    .Q(\rbzero.wall_tracer.trackDistY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _20972_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00561_),
    .Q(\rbzero.wall_tracer.trackDistY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _20973_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00562_),
    .Q(\rbzero.wall_tracer.trackDistY[1] ));
 sky130_fd_sc_hd__dfxtp_1 _20974_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00563_),
    .Q(\rbzero.wall_tracer.trackDistY[2] ));
 sky130_fd_sc_hd__dfxtp_1 _20975_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00564_),
    .Q(\rbzero.wall_tracer.trackDistY[3] ));
 sky130_fd_sc_hd__dfxtp_1 _20976_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00565_),
    .Q(\rbzero.wall_tracer.trackDistY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _20977_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00566_),
    .Q(\rbzero.wall_tracer.trackDistY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _20978_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00567_),
    .Q(\rbzero.wall_tracer.trackDistY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _20979_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00568_),
    .Q(\rbzero.wall_tracer.trackDistY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _20980_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00569_),
    .Q(\rbzero.wall_tracer.trackDistY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _20981_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00570_),
    .Q(\rbzero.wall_tracer.trackDistY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _20982_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00571_),
    .Q(\rbzero.wall_tracer.trackDistY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _20983_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00572_),
    .Q(\rbzero.spi_registers.new_texadd[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _20984_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00573_),
    .Q(\rbzero.spi_registers.new_texadd[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _20985_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00574_),
    .Q(\rbzero.spi_registers.new_texadd[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _20986_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00575_),
    .Q(\rbzero.spi_registers.new_texadd[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _20987_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00576_),
    .Q(\rbzero.spi_registers.new_texadd[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _20988_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00577_),
    .Q(\rbzero.spi_registers.new_texadd[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _20989_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00578_),
    .Q(\rbzero.spi_registers.new_texadd[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _20990_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00579_),
    .Q(\rbzero.spi_registers.new_texadd[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _20991_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00580_),
    .Q(\rbzero.spi_registers.new_texadd[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _20992_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00581_),
    .Q(\rbzero.spi_registers.new_texadd[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _20993_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00582_),
    .Q(\rbzero.spi_registers.new_texadd[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _20994_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00583_),
    .Q(\rbzero.spi_registers.new_texadd[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _20995_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00584_),
    .Q(\rbzero.spi_registers.new_texadd[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _20996_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00585_),
    .Q(\rbzero.spi_registers.new_texadd[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _20997_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00586_),
    .Q(\rbzero.spi_registers.new_texadd[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _20998_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00587_),
    .Q(\rbzero.spi_registers.new_texadd[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _20999_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00588_),
    .Q(\rbzero.spi_registers.new_texadd[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21000_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00589_),
    .Q(\rbzero.spi_registers.new_texadd[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21001_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00590_),
    .Q(\rbzero.spi_registers.new_texadd[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21002_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00591_),
    .Q(\rbzero.spi_registers.new_texadd[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21003_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00592_),
    .Q(\rbzero.spi_registers.new_texadd[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21004_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00593_),
    .Q(\rbzero.spi_registers.new_texadd[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21005_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00594_),
    .Q(\rbzero.spi_registers.new_texadd[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21006_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00595_),
    .Q(\rbzero.spi_registers.new_texadd[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21007_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00596_),
    .Q(\rbzero.wall_tracer.rayAddendX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21008_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00597_),
    .Q(\rbzero.wall_tracer.rayAddendX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21009_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00598_),
    .Q(\rbzero.wall_tracer.rayAddendX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21010_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00599_),
    .Q(\rbzero.wall_tracer.rayAddendX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21011_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00600_),
    .Q(\rbzero.wall_tracer.rayAddendX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21012_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00601_),
    .Q(\rbzero.wall_tracer.rayAddendX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21013_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00602_),
    .Q(\rbzero.wall_tracer.rayAddendX[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21014_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00603_),
    .Q(\rbzero.wall_tracer.rayAddendX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21015_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00604_),
    .Q(\rbzero.wall_tracer.rayAddendX[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21016_ (.CLK(clknet_3_5_0_i_clk),
    .D(_00605_),
    .Q(\rbzero.wall_tracer.rayAddendX[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21017_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00606_),
    .Q(\rbzero.wall_tracer.rayAddendX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21018_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00607_),
    .Q(\rbzero.wall_tracer.rayAddendX[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21019_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00608_),
    .Q(\rbzero.wall_tracer.rayAddendX[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21020_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00609_),
    .Q(\rbzero.wall_tracer.rayAddendX[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21021_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00610_),
    .Q(\rbzero.wall_tracer.rayAddendX[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21022_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00611_),
    .Q(\rbzero.wall_tracer.rayAddendX[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21023_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00612_),
    .Q(\rbzero.map_rom.d6 ));
 sky130_fd_sc_hd__dfxtp_2 _21024_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00613_),
    .Q(\rbzero.map_rom.c6 ));
 sky130_fd_sc_hd__dfxtp_2 _21025_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00614_),
    .Q(\rbzero.map_rom.b6 ));
 sky130_fd_sc_hd__dfxtp_2 _21026_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00615_),
    .Q(\rbzero.map_rom.a6 ));
 sky130_fd_sc_hd__dfxtp_4 _21027_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00616_),
    .Q(\rbzero.map_rom.i_row[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21028_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00617_),
    .Q(\rbzero.wall_tracer.mapY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21029_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00618_),
    .Q(\rbzero.map_rom.f4 ));
 sky130_fd_sc_hd__dfxtp_1 _21030_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00619_),
    .Q(\rbzero.map_rom.f3 ));
 sky130_fd_sc_hd__dfxtp_2 _21031_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00620_),
    .Q(\rbzero.map_rom.f2 ));
 sky130_fd_sc_hd__dfxtp_2 _21032_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00621_),
    .Q(\rbzero.map_rom.f1 ));
 sky130_fd_sc_hd__dfxtp_2 _21033_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00622_),
    .Q(\rbzero.map_rom.i_col[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21034_ (.CLK(clknet_leaf_46_i_clk),
    .D(_00623_),
    .Q(\rbzero.wall_tracer.mapX[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21035_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00624_),
    .Q(\rbzero.wall_tracer.rayAddendY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21036_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00625_),
    .Q(\rbzero.wall_tracer.rayAddendY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21037_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00626_),
    .Q(\rbzero.wall_tracer.rayAddendY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21038_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00627_),
    .Q(\rbzero.wall_tracer.rayAddendY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21039_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00628_),
    .Q(\rbzero.wall_tracer.rayAddendY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21040_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00629_),
    .Q(\rbzero.wall_tracer.rayAddendY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21041_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00630_),
    .Q(\rbzero.wall_tracer.rayAddendY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21042_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00631_),
    .Q(\rbzero.wall_tracer.rayAddendY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21043_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00632_),
    .Q(\rbzero.wall_tracer.rayAddendY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21044_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00633_),
    .Q(\rbzero.wall_tracer.rayAddendY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21045_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00634_),
    .Q(\rbzero.wall_tracer.rayAddendY[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21046_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00635_),
    .Q(\rbzero.wall_tracer.rayAddendY[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21047_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00636_),
    .Q(\rbzero.wall_tracer.rayAddendY[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21048_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00637_),
    .Q(\rbzero.wall_tracer.rayAddendY[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21049_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00638_),
    .Q(\rbzero.wall_tracer.rayAddendY[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21050_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00639_),
    .Q(\rbzero.wall_tracer.rayAddendY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21051_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00640_),
    .Q(\rbzero.spi_registers.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21052_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00641_),
    .Q(\rbzero.spi_registers.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21053_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00642_),
    .Q(\rbzero.spi_registers.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21054_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00643_),
    .Q(\rbzero.spi_registers.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21055_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00644_),
    .Q(\rbzero.spi_registers.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21056_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00645_),
    .Q(\rbzero.spi_registers.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21057_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00646_),
    .Q(\rbzero.spi_registers.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21058_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00647_),
    .Q(\rbzero.pov.ready_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21059_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00648_),
    .Q(\rbzero.pov.ready_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21060_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00649_),
    .Q(\rbzero.pov.ready_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21061_ (.CLK(clknet_leaf_98_i_clk),
    .D(_00650_),
    .Q(\rbzero.pov.ready_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21062_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00651_),
    .Q(\rbzero.pov.ready_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21063_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00652_),
    .Q(\rbzero.pov.ready_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21064_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00653_),
    .Q(\rbzero.pov.ready_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21065_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00654_),
    .Q(\rbzero.pov.ready_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21066_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00655_),
    .Q(\rbzero.pov.ready_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21067_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00656_),
    .Q(\rbzero.pov.ready_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21068_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00657_),
    .Q(\rbzero.pov.ready_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21069_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00658_),
    .Q(\rbzero.pov.ready_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21070_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00659_),
    .Q(\rbzero.pov.ready_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21071_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00660_),
    .Q(\rbzero.pov.ready_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21072_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00661_),
    .Q(\rbzero.pov.ready_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21073_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00662_),
    .Q(\rbzero.pov.ready_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21074_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00663_),
    .Q(\rbzero.pov.ready_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21075_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00664_),
    .Q(\rbzero.pov.ready_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21076_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00665_),
    .Q(\rbzero.pov.ready_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21077_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00666_),
    .Q(\rbzero.pov.ready_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21078_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00667_),
    .Q(\rbzero.pov.ready_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21079_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00668_),
    .Q(\rbzero.pov.ready_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21080_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00669_),
    .Q(\rbzero.pov.ready_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21081_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00670_),
    .Q(\rbzero.pov.ready_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21082_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00671_),
    .Q(\rbzero.pov.ready_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21083_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00672_),
    .Q(\rbzero.pov.ready_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21084_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00673_),
    .Q(\rbzero.pov.ready_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21085_ (.CLK(clknet_leaf_88_i_clk),
    .D(_00674_),
    .Q(\rbzero.pov.ready_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21086_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00675_),
    .Q(\rbzero.pov.ready_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21087_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00676_),
    .Q(\rbzero.pov.ready_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21088_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00677_),
    .Q(\rbzero.pov.ready_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21089_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00678_),
    .Q(\rbzero.pov.ready_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21090_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00679_),
    .Q(\rbzero.pov.ready_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21091_ (.CLK(clknet_leaf_97_i_clk),
    .D(_00680_),
    .Q(\rbzero.pov.ready_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21092_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00681_),
    .Q(\rbzero.pov.ready_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21093_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00682_),
    .Q(\rbzero.pov.ready_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21094_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00683_),
    .Q(\rbzero.pov.ready_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21095_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00684_),
    .Q(\rbzero.pov.ready_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21096_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00685_),
    .Q(\rbzero.pov.ready_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21097_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00686_),
    .Q(\rbzero.pov.ready_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21098_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00687_),
    .Q(\rbzero.pov.ready_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21099_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00688_),
    .Q(\rbzero.pov.ready_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21100_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00689_),
    .Q(\rbzero.pov.ready_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21101_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00690_),
    .Q(\rbzero.pov.ready_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21102_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00691_),
    .Q(\rbzero.pov.ready_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21103_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00692_),
    .Q(\rbzero.pov.ready_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21104_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00693_),
    .Q(\rbzero.pov.ready_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21105_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00694_),
    .Q(\rbzero.pov.ready_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21106_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00695_),
    .Q(\rbzero.pov.ready_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21107_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00696_),
    .Q(\rbzero.pov.ready_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21108_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00697_),
    .Q(\rbzero.pov.ready_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21109_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00698_),
    .Q(\rbzero.pov.ready_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21110_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00699_),
    .Q(\rbzero.pov.ready_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21111_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00700_),
    .Q(\rbzero.pov.ready_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21112_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00701_),
    .Q(\rbzero.pov.ready_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21113_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00702_),
    .Q(\rbzero.pov.ready_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21114_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00703_),
    .Q(\rbzero.pov.ready_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21115_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00704_),
    .Q(\rbzero.pov.ready_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21116_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00705_),
    .Q(\rbzero.pov.ready_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21117_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00706_),
    .Q(\rbzero.pov.ready_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21118_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00707_),
    .Q(\rbzero.pov.ready_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21119_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00708_),
    .Q(\rbzero.pov.ready_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21120_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00709_),
    .Q(\rbzero.pov.ready_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21121_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00710_),
    .Q(\rbzero.pov.ready_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21122_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00711_),
    .Q(\rbzero.pov.ready_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21123_ (.CLK(clknet_leaf_91_i_clk),
    .D(_00712_),
    .Q(\rbzero.pov.ready_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21124_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00713_),
    .Q(\rbzero.pov.ready_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21125_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00714_),
    .Q(\rbzero.pov.ready_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21126_ (.CLK(clknet_leaf_92_i_clk),
    .D(_00715_),
    .Q(\rbzero.pov.ready_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21127_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00716_),
    .Q(\rbzero.pov.ready_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21128_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00717_),
    .Q(\rbzero.pov.ready_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21129_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00718_),
    .Q(\rbzero.pov.ready_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21130_ (.CLK(clknet_leaf_93_i_clk),
    .D(_00719_),
    .Q(\rbzero.pov.ready_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21131_ (.CLK(clknet_leaf_96_i_clk),
    .D(_00720_),
    .Q(\rbzero.pov.ready_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21132_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00721_),
    .Q(\rbzero.spi_registers.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21133_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00722_),
    .Q(\rbzero.spi_registers.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21134_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00723_),
    .Q(\rbzero.spi_registers.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21135_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00724_),
    .Q(\rbzero.spi_registers.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21136_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00725_),
    .Q(\rbzero.spi_registers.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21137_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00726_),
    .Q(\rbzero.spi_registers.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21138_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00727_),
    .Q(\rbzero.spi_registers.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21139_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00728_),
    .Q(\rbzero.spi_registers.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_2 _21140_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00729_),
    .Q(\rbzero.spi_registers.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_2 _21141_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00730_),
    .Q(\rbzero.spi_registers.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_2 _21142_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00731_),
    .Q(\rbzero.spi_registers.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21143_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00732_),
    .Q(\rbzero.spi_registers.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_2 _21144_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00733_),
    .Q(\rbzero.spi_registers.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_2 _21145_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00734_),
    .Q(\rbzero.spi_registers.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_2 _21146_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00735_),
    .Q(\rbzero.spi_registers.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_2 _21147_ (.CLK(clknet_leaf_99_i_clk),
    .D(_00736_),
    .Q(\rbzero.spi_registers.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21148_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00737_),
    .Q(\rbzero.spi_registers.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21149_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00738_),
    .Q(\rbzero.spi_registers.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21150_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00739_),
    .Q(\rbzero.spi_registers.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_2 _21151_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00740_),
    .Q(\rbzero.spi_registers.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21152_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00741_),
    .Q(\rbzero.spi_registers.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21153_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00742_),
    .Q(\rbzero.spi_registers.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21154_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00743_),
    .Q(\rbzero.spi_registers.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21155_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00744_),
    .Q(\rbzero.spi_registers.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21156_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00745_),
    .Q(\rbzero.spi_registers.spi_cmd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21157_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00746_),
    .Q(\rbzero.spi_registers.spi_cmd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21158_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00747_),
    .Q(\rbzero.spi_registers.spi_cmd[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21159_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00748_),
    .Q(\rbzero.spi_registers.spi_cmd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21160_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00749_),
    .Q(\rbzero.spi_registers.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21161_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00750_),
    .Q(\rbzero.spi_registers.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21162_ (.CLK(clknet_leaf_94_i_clk),
    .D(_00751_),
    .Q(\rbzero.spi_registers.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21163_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00752_),
    .Q(\rbzero.spi_registers.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21164_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00753_),
    .Q(\rbzero.spi_registers.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21165_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00754_),
    .Q(\rbzero.spi_registers.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21166_ (.CLK(clknet_leaf_95_i_clk),
    .D(_00755_),
    .Q(\rbzero.spi_registers.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21167_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00756_),
    .Q(\rbzero.map_overlay.i_otherx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21168_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00757_),
    .Q(\rbzero.map_overlay.i_otherx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21169_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00758_),
    .Q(\rbzero.map_overlay.i_otherx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21170_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00759_),
    .Q(\rbzero.map_overlay.i_otherx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21171_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00760_),
    .Q(\rbzero.map_overlay.i_otherx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21172_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00761_),
    .Q(\rbzero.map_overlay.i_othery[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21173_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00762_),
    .Q(\rbzero.map_overlay.i_othery[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21174_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00763_),
    .Q(\rbzero.map_overlay.i_othery[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21175_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00764_),
    .Q(\rbzero.map_overlay.i_othery[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21176_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00765_),
    .Q(\rbzero.map_overlay.i_othery[4] ));
 sky130_fd_sc_hd__dfxtp_2 _21177_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00766_),
    .Q(\rbzero.row_render.vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21178_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00767_),
    .Q(\rbzero.map_overlay.i_mapdx[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21179_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00768_),
    .Q(\rbzero.map_overlay.i_mapdx[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21180_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00769_),
    .Q(\rbzero.map_overlay.i_mapdx[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21181_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00770_),
    .Q(\rbzero.map_overlay.i_mapdx[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21182_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00771_),
    .Q(\rbzero.map_overlay.i_mapdx[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21183_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00772_),
    .Q(\rbzero.map_overlay.i_mapdx[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21184_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00773_),
    .Q(\rbzero.map_overlay.i_mapdy[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21185_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00774_),
    .Q(\rbzero.map_overlay.i_mapdy[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21186_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00775_),
    .Q(\rbzero.map_overlay.i_mapdy[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21187_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00776_),
    .Q(\rbzero.map_overlay.i_mapdy[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21188_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00777_),
    .Q(\rbzero.map_overlay.i_mapdy[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21189_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00778_),
    .Q(\rbzero.map_overlay.i_mapdy[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21190_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00779_),
    .Q(\rbzero.mapdxw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21191_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00780_),
    .Q(\rbzero.mapdxw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21192_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00781_),
    .Q(\rbzero.mapdyw[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21193_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00782_),
    .Q(\rbzero.mapdyw[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21194_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00783_),
    .Q(\rbzero.spi_registers.texadd0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21195_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00784_),
    .Q(\rbzero.spi_registers.texadd0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21196_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00785_),
    .Q(\rbzero.spi_registers.texadd0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21197_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00786_),
    .Q(\rbzero.spi_registers.texadd0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21198_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00787_),
    .Q(\rbzero.spi_registers.texadd0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21199_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00788_),
    .Q(\rbzero.spi_registers.texadd0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21200_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00789_),
    .Q(\rbzero.spi_registers.texadd0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21201_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00790_),
    .Q(\rbzero.spi_registers.texadd0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21202_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00791_),
    .Q(\rbzero.spi_registers.texadd0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21203_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00792_),
    .Q(\rbzero.spi_registers.texadd0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21204_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00793_),
    .Q(\rbzero.spi_registers.texadd0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21205_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00794_),
    .Q(\rbzero.spi_registers.texadd0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21206_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00795_),
    .Q(\rbzero.spi_registers.texadd0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21207_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00796_),
    .Q(\rbzero.spi_registers.texadd0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21208_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00797_),
    .Q(\rbzero.spi_registers.texadd0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21209_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00798_),
    .Q(\rbzero.spi_registers.texadd0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21210_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00799_),
    .Q(\rbzero.spi_registers.texadd0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21211_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00800_),
    .Q(\rbzero.spi_registers.texadd0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21212_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00801_),
    .Q(\rbzero.spi_registers.texadd0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21213_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00802_),
    .Q(\rbzero.spi_registers.texadd0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21214_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00803_),
    .Q(\rbzero.spi_registers.texadd0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21215_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00804_),
    .Q(\rbzero.spi_registers.texadd0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21216_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00805_),
    .Q(\rbzero.spi_registers.texadd0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21217_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00806_),
    .Q(\rbzero.spi_registers.texadd0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21218_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00807_),
    .Q(\rbzero.spi_registers.texadd1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21219_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00808_),
    .Q(\rbzero.spi_registers.texadd1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21220_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00809_),
    .Q(\rbzero.spi_registers.texadd1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21221_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00810_),
    .Q(\rbzero.spi_registers.texadd1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21222_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00811_),
    .Q(\rbzero.spi_registers.texadd1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21223_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00812_),
    .Q(\rbzero.spi_registers.texadd1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21224_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00813_),
    .Q(\rbzero.spi_registers.texadd1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21225_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00814_),
    .Q(\rbzero.spi_registers.texadd1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21226_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00815_),
    .Q(\rbzero.spi_registers.texadd1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21227_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00816_),
    .Q(\rbzero.spi_registers.texadd1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21228_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00817_),
    .Q(\rbzero.spi_registers.texadd1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21229_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00818_),
    .Q(\rbzero.spi_registers.texadd1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21230_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00819_),
    .Q(\rbzero.spi_registers.texadd1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21231_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00820_),
    .Q(\rbzero.spi_registers.texadd1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21232_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00821_),
    .Q(\rbzero.spi_registers.texadd1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21233_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00822_),
    .Q(\rbzero.spi_registers.texadd1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21234_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00823_),
    .Q(\rbzero.spi_registers.texadd1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21235_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00824_),
    .Q(\rbzero.spi_registers.texadd1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21236_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00825_),
    .Q(\rbzero.spi_registers.texadd1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21237_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00826_),
    .Q(\rbzero.spi_registers.texadd1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21238_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00827_),
    .Q(\rbzero.spi_registers.texadd1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21239_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00828_),
    .Q(\rbzero.spi_registers.texadd1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21240_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00829_),
    .Q(\rbzero.spi_registers.texadd1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21241_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00830_),
    .Q(\rbzero.spi_registers.texadd1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21242_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00831_),
    .Q(\rbzero.spi_registers.texadd2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21243_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00832_),
    .Q(\rbzero.spi_registers.texadd2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21244_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00833_),
    .Q(\rbzero.spi_registers.texadd2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21245_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00834_),
    .Q(\rbzero.spi_registers.texadd2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21246_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00835_),
    .Q(\rbzero.spi_registers.texadd2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21247_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00836_),
    .Q(\rbzero.spi_registers.texadd2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21248_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00837_),
    .Q(\rbzero.spi_registers.texadd2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21249_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00838_),
    .Q(\rbzero.spi_registers.texadd2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21250_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00839_),
    .Q(\rbzero.spi_registers.texadd2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21251_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00840_),
    .Q(\rbzero.spi_registers.texadd2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21252_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00841_),
    .Q(\rbzero.spi_registers.texadd2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21253_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00842_),
    .Q(\rbzero.spi_registers.texadd2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21254_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00843_),
    .Q(\rbzero.spi_registers.texadd2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21255_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00844_),
    .Q(\rbzero.spi_registers.texadd2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21256_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00845_),
    .Q(\rbzero.spi_registers.texadd2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21257_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00846_),
    .Q(\rbzero.spi_registers.texadd2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21258_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00847_),
    .Q(\rbzero.spi_registers.texadd2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21259_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00848_),
    .Q(\rbzero.spi_registers.texadd2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21260_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00849_),
    .Q(\rbzero.spi_registers.texadd2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21261_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00850_),
    .Q(\rbzero.spi_registers.texadd2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21262_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00851_),
    .Q(\rbzero.spi_registers.texadd2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21263_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00852_),
    .Q(\rbzero.spi_registers.texadd2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21264_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00853_),
    .Q(\rbzero.spi_registers.texadd2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21265_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00854_),
    .Q(\rbzero.spi_registers.texadd2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21266_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00855_),
    .Q(\rbzero.spi_registers.texadd3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21267_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00856_),
    .Q(\rbzero.spi_registers.texadd3[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21268_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00857_),
    .Q(\rbzero.spi_registers.texadd3[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21269_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00858_),
    .Q(\rbzero.spi_registers.texadd3[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21270_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00859_),
    .Q(\rbzero.spi_registers.texadd3[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21271_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00860_),
    .Q(\rbzero.spi_registers.texadd3[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21272_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00861_),
    .Q(\rbzero.spi_registers.texadd3[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21273_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00862_),
    .Q(\rbzero.spi_registers.texadd3[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21274_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00863_),
    .Q(\rbzero.spi_registers.texadd3[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21275_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00864_),
    .Q(\rbzero.spi_registers.texadd3[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21276_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00865_),
    .Q(\rbzero.spi_registers.texadd3[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21277_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00866_),
    .Q(\rbzero.spi_registers.texadd3[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21278_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00867_),
    .Q(\rbzero.spi_registers.texadd3[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21279_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00868_),
    .Q(\rbzero.spi_registers.texadd3[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21280_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00869_),
    .Q(\rbzero.spi_registers.texadd3[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21281_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00870_),
    .Q(\rbzero.spi_registers.texadd3[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21282_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00871_),
    .Q(\rbzero.spi_registers.texadd3[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21283_ (.CLK(clknet_leaf_100_i_clk),
    .D(_00872_),
    .Q(\rbzero.spi_registers.texadd3[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21284_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00873_),
    .Q(\rbzero.spi_registers.texadd3[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21285_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00874_),
    .Q(\rbzero.spi_registers.texadd3[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21286_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00875_),
    .Q(\rbzero.spi_registers.texadd3[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21287_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00876_),
    .Q(\rbzero.spi_registers.texadd3[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21288_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00877_),
    .Q(\rbzero.spi_registers.texadd3[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21289_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00878_),
    .Q(\rbzero.spi_registers.texadd3[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21290_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00879_),
    .Q(\rbzero.floor_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21291_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00880_),
    .Q(\rbzero.floor_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21292_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00881_),
    .Q(\rbzero.floor_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21293_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00882_),
    .Q(\rbzero.floor_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21294_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00883_),
    .Q(\rbzero.floor_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21295_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00884_),
    .Q(\rbzero.floor_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21296_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00885_),
    .Q(\rbzero.color_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21297_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00886_),
    .Q(\rbzero.color_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21298_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00887_),
    .Q(\rbzero.color_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21299_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00888_),
    .Q(\rbzero.color_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21300_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00889_),
    .Q(\rbzero.color_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21301_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00890_),
    .Q(\rbzero.color_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21302_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00891_),
    .Q(\rbzero.color_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21303_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00892_),
    .Q(\rbzero.color_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21304_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00893_),
    .Q(\rbzero.color_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21305_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00894_),
    .Q(\rbzero.color_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21306_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00895_),
    .Q(\rbzero.color_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21307_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00896_),
    .Q(\rbzero.color_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21308_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00897_),
    .Q(\rbzero.spi_registers.vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21309_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00898_),
    .Q(\rbzero.spi_registers.vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21310_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00899_),
    .Q(\rbzero.spi_registers.vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21311_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00900_),
    .Q(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21312_ (.CLK(clknet_leaf_34_i_clk),
    .D(_00901_),
    .Q(\rbzero.spi_registers.vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21313_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00902_),
    .Q(\rbzero.spi_registers.vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21314_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00903_),
    .Q(\rbzero.spi_registers.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21315_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00904_),
    .Q(\rbzero.spi_registers.new_sky[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21316_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00905_),
    .Q(\rbzero.spi_registers.new_sky[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21317_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00906_),
    .Q(\rbzero.spi_registers.new_sky[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21318_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00907_),
    .Q(\rbzero.spi_registers.new_sky[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21319_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00908_),
    .Q(\rbzero.spi_registers.new_sky[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21320_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00909_),
    .Q(\rbzero.spi_registers.new_sky[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21321_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00910_),
    .Q(\rbzero.spi_registers.got_new_sky ));
 sky130_fd_sc_hd__dfxtp_1 _21322_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00911_),
    .Q(\rbzero.spi_registers.new_floor[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21323_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00912_),
    .Q(\rbzero.spi_registers.new_floor[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21324_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00913_),
    .Q(\rbzero.spi_registers.new_floor[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21325_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00914_),
    .Q(\rbzero.spi_registers.new_floor[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21326_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00915_),
    .Q(\rbzero.spi_registers.new_floor[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21327_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00916_),
    .Q(\rbzero.spi_registers.new_floor[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21328_ (.CLK(clknet_leaf_30_i_clk),
    .D(_00917_),
    .Q(\rbzero.spi_registers.got_new_floor ));
 sky130_fd_sc_hd__dfxtp_1 _21329_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00918_),
    .Q(\rbzero.spi_registers.new_leak[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21330_ (.CLK(clknet_leaf_33_i_clk),
    .D(_00919_),
    .Q(\rbzero.spi_registers.new_leak[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21331_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00920_),
    .Q(\rbzero.spi_registers.new_leak[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21332_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00921_),
    .Q(\rbzero.spi_registers.new_leak[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21333_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00922_),
    .Q(\rbzero.spi_registers.new_leak[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21334_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00923_),
    .Q(\rbzero.spi_registers.new_leak[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21335_ (.CLK(clknet_leaf_31_i_clk),
    .D(_00924_),
    .Q(\rbzero.spi_registers.got_new_leak ));
 sky130_fd_sc_hd__dfxtp_1 _21336_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00925_),
    .Q(\rbzero.spi_registers.new_other[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21337_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00926_),
    .Q(\rbzero.spi_registers.new_other[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21338_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00927_),
    .Q(\rbzero.spi_registers.new_other[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21339_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00928_),
    .Q(\rbzero.spi_registers.new_other[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21340_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00929_),
    .Q(\rbzero.spi_registers.new_other[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21341_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00930_),
    .Q(\rbzero.spi_registers.new_other[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21342_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00931_),
    .Q(\rbzero.spi_registers.new_other[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21343_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00932_),
    .Q(\rbzero.spi_registers.new_other[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21344_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00933_),
    .Q(\rbzero.spi_registers.new_other[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21345_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00934_),
    .Q(\rbzero.spi_registers.new_other[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21346_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00935_),
    .Q(\rbzero.spi_registers.got_new_other ));
 sky130_fd_sc_hd__dfxtp_1 _21347_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00936_),
    .Q(\rbzero.spi_registers.new_vshift[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21348_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00937_),
    .Q(\rbzero.spi_registers.new_vshift[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21349_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00938_),
    .Q(\rbzero.spi_registers.new_vshift[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21350_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00939_),
    .Q(\rbzero.spi_registers.new_vshift[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21351_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00940_),
    .Q(\rbzero.spi_registers.new_vshift[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21352_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00941_),
    .Q(\rbzero.spi_registers.new_vshift[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21353_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00942_),
    .Q(\rbzero.spi_registers.got_new_vshift ));
 sky130_fd_sc_hd__dfxtp_1 _21354_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00943_),
    .Q(\rbzero.spi_registers.new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21355_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00944_),
    .Q(\rbzero.spi_registers.got_new_vinf ));
 sky130_fd_sc_hd__dfxtp_1 _21356_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00945_),
    .Q(\rbzero.spi_registers.new_mapd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21357_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00946_),
    .Q(\rbzero.spi_registers.new_mapd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21358_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00947_),
    .Q(\rbzero.spi_registers.new_mapd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21359_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00948_),
    .Q(\rbzero.spi_registers.new_mapd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21360_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00949_),
    .Q(\rbzero.spi_registers.new_mapd[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21361_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00950_),
    .Q(\rbzero.spi_registers.new_mapd[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21362_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00951_),
    .Q(\rbzero.spi_registers.new_mapd[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21363_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00952_),
    .Q(\rbzero.spi_registers.new_mapd[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21364_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00953_),
    .Q(\rbzero.spi_registers.new_mapd[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21365_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00954_),
    .Q(\rbzero.spi_registers.new_mapd[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21366_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00955_),
    .Q(\rbzero.spi_registers.new_mapd[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21367_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00956_),
    .Q(\rbzero.spi_registers.new_mapd[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21368_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00957_),
    .Q(\rbzero.spi_registers.new_mapd[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21369_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00958_),
    .Q(\rbzero.spi_registers.new_mapd[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21370_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00959_),
    .Q(\rbzero.spi_registers.new_mapd[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21371_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00960_),
    .Q(\rbzero.spi_registers.new_mapd[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21372_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00961_),
    .Q(\rbzero.spi_registers.got_new_mapd ));
 sky130_fd_sc_hd__dfxtp_1 _21373_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00962_),
    .Q(\rbzero.spi_registers.got_new_texadd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21374_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00963_),
    .Q(\rbzero.spi_registers.got_new_texadd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21375_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00964_),
    .Q(\rbzero.spi_registers.got_new_texadd[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21376_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00965_),
    .Q(\rbzero.spi_registers.got_new_texadd[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21377_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00966_),
    .Q(\rbzero.spi_registers.new_texadd[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21378_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00967_),
    .Q(\rbzero.spi_registers.new_texadd[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21379_ (.CLK(clknet_leaf_29_i_clk),
    .D(_00968_),
    .Q(\rbzero.spi_registers.new_texadd[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21380_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00969_),
    .Q(\rbzero.spi_registers.new_texadd[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21381_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00970_),
    .Q(\rbzero.spi_registers.new_texadd[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21382_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00971_),
    .Q(\rbzero.spi_registers.new_texadd[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21383_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00972_),
    .Q(\rbzero.spi_registers.new_texadd[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21384_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00973_),
    .Q(\rbzero.spi_registers.new_texadd[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21385_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00974_),
    .Q(\rbzero.spi_registers.new_texadd[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21386_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00975_),
    .Q(\rbzero.spi_registers.new_texadd[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21387_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00976_),
    .Q(\rbzero.spi_registers.new_texadd[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21388_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00977_),
    .Q(\rbzero.spi_registers.new_texadd[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21389_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00978_),
    .Q(\rbzero.spi_registers.new_texadd[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21390_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00979_),
    .Q(\rbzero.spi_registers.new_texadd[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21391_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00980_),
    .Q(\rbzero.spi_registers.new_texadd[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21392_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00981_),
    .Q(\rbzero.spi_registers.new_texadd[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21393_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00982_),
    .Q(\rbzero.spi_registers.new_texadd[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21394_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00983_),
    .Q(\rbzero.spi_registers.new_texadd[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21395_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00984_),
    .Q(\rbzero.spi_registers.new_texadd[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21396_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00985_),
    .Q(\rbzero.spi_registers.new_texadd[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21397_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00986_),
    .Q(\rbzero.spi_registers.new_texadd[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21398_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00987_),
    .Q(\rbzero.spi_registers.new_texadd[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21399_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00988_),
    .Q(\rbzero.spi_registers.new_texadd[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21400_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00989_),
    .Q(\rbzero.spi_registers.new_texadd[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21401_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00990_),
    .Q(\rbzero.spi_registers.new_texadd[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21402_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00991_),
    .Q(\rbzero.spi_registers.new_texadd[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21403_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00992_),
    .Q(\rbzero.spi_registers.new_texadd[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21404_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00993_),
    .Q(\rbzero.spi_registers.new_texadd[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21405_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00994_),
    .Q(\rbzero.spi_registers.new_texadd[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21406_ (.CLK(clknet_leaf_28_i_clk),
    .D(_00995_),
    .Q(\rbzero.spi_registers.new_texadd[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21407_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00996_),
    .Q(\rbzero.spi_registers.new_texadd[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21408_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00997_),
    .Q(\rbzero.spi_registers.new_texadd[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21409_ (.CLK(clknet_leaf_24_i_clk),
    .D(_00998_),
    .Q(\rbzero.spi_registers.new_texadd[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21410_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00999_),
    .Q(\rbzero.spi_registers.new_texadd[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21411_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01000_),
    .Q(\rbzero.spi_registers.new_texadd[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21412_ (.CLK(clknet_leaf_2_i_clk),
    .D(_01001_),
    .Q(\rbzero.spi_registers.new_texadd[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21413_ (.CLK(clknet_leaf_12_i_clk),
    .D(_01002_),
    .Q(\rbzero.spi_registers.new_texadd[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21414_ (.CLK(clknet_leaf_1_i_clk),
    .D(_01003_),
    .Q(\rbzero.spi_registers.new_texadd[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21415_ (.CLK(clknet_leaf_11_i_clk),
    .D(_01004_),
    .Q(\rbzero.spi_registers.new_texadd[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21416_ (.CLK(clknet_leaf_1_i_clk),
    .D(_01005_),
    .Q(\rbzero.spi_registers.new_texadd[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21417_ (.CLK(clknet_leaf_2_i_clk),
    .D(_01006_),
    .Q(\rbzero.spi_registers.new_texadd[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21418_ (.CLK(clknet_leaf_2_i_clk),
    .D(_01007_),
    .Q(\rbzero.spi_registers.new_texadd[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21419_ (.CLK(clknet_leaf_4_i_clk),
    .D(_01008_),
    .Q(\rbzero.spi_registers.new_texadd[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21420_ (.CLK(clknet_leaf_4_i_clk),
    .D(_01009_),
    .Q(\rbzero.spi_registers.new_texadd[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21421_ (.CLK(clknet_leaf_4_i_clk),
    .D(_01010_),
    .Q(\rbzero.spi_registers.new_texadd[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21422_ (.CLK(clknet_leaf_4_i_clk),
    .D(_01011_),
    .Q(\rbzero.spi_registers.new_texadd[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21423_ (.CLK(clknet_leaf_25_i_clk),
    .D(_01012_),
    .Q(\rbzero.spi_registers.new_texadd[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21424_ (.CLK(clknet_leaf_6_i_clk),
    .D(_01013_),
    .Q(\rbzero.spi_registers.new_texadd[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21425_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01014_),
    .Q(\rbzero.pov.ready ));
 sky130_fd_sc_hd__dfxtp_1 _21426_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01015_),
    .Q(\rbzero.pov.spi_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21427_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01016_),
    .Q(\rbzero.pov.spi_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21428_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01017_),
    .Q(\rbzero.pov.spi_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21429_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01018_),
    .Q(\rbzero.pov.spi_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21430_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01019_),
    .Q(\rbzero.pov.spi_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21431_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01020_),
    .Q(\rbzero.pov.spi_counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21432_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01021_),
    .Q(\rbzero.pov.spi_counter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21433_ (.CLK(net151),
    .D(_01022_),
    .Q(\rbzero.tex_b0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21434_ (.CLK(net152),
    .D(_01023_),
    .Q(\rbzero.tex_b0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21435_ (.CLK(net153),
    .D(_01024_),
    .Q(\rbzero.tex_b0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21436_ (.CLK(net154),
    .D(_01025_),
    .Q(\rbzero.tex_b0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21437_ (.CLK(net155),
    .D(_01026_),
    .Q(\rbzero.tex_b0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21438_ (.CLK(net156),
    .D(_01027_),
    .Q(\rbzero.tex_b0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21439_ (.CLK(net157),
    .D(_01028_),
    .Q(\rbzero.tex_b0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21440_ (.CLK(net158),
    .D(_01029_),
    .Q(\rbzero.tex_b0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21441_ (.CLK(net159),
    .D(_01030_),
    .Q(\rbzero.tex_b0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21442_ (.CLK(net160),
    .D(_01031_),
    .Q(\rbzero.tex_b0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21443_ (.CLK(net161),
    .D(_01032_),
    .Q(\rbzero.tex_b0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21444_ (.CLK(net162),
    .D(_01033_),
    .Q(\rbzero.tex_b0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21445_ (.CLK(net163),
    .D(_01034_),
    .Q(\rbzero.tex_b0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21446_ (.CLK(net164),
    .D(_01035_),
    .Q(\rbzero.tex_b0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21447_ (.CLK(net165),
    .D(_01036_),
    .Q(\rbzero.tex_b0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21448_ (.CLK(net166),
    .D(_01037_),
    .Q(\rbzero.tex_b0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21449_ (.CLK(net167),
    .D(_01038_),
    .Q(\rbzero.tex_b0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21450_ (.CLK(net168),
    .D(_01039_),
    .Q(\rbzero.tex_b0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21451_ (.CLK(net169),
    .D(_01040_),
    .Q(\rbzero.tex_b0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21452_ (.CLK(net170),
    .D(_01041_),
    .Q(\rbzero.tex_b0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21453_ (.CLK(net171),
    .D(_01042_),
    .Q(\rbzero.tex_b0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21454_ (.CLK(net172),
    .D(_01043_),
    .Q(\rbzero.tex_b0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21455_ (.CLK(net173),
    .D(_01044_),
    .Q(\rbzero.tex_b0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21456_ (.CLK(net174),
    .D(_01045_),
    .Q(\rbzero.tex_b0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21457_ (.CLK(net175),
    .D(_01046_),
    .Q(\rbzero.tex_b0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21458_ (.CLK(net176),
    .D(_01047_),
    .Q(\rbzero.tex_b0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21459_ (.CLK(net177),
    .D(_01048_),
    .Q(\rbzero.tex_b0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21460_ (.CLK(net178),
    .D(_01049_),
    .Q(\rbzero.tex_b0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21461_ (.CLK(net179),
    .D(_01050_),
    .Q(\rbzero.tex_b0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21462_ (.CLK(net180),
    .D(_01051_),
    .Q(\rbzero.tex_b0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21463_ (.CLK(net181),
    .D(_01052_),
    .Q(\rbzero.tex_b0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21464_ (.CLK(net182),
    .D(_01053_),
    .Q(\rbzero.tex_b0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21465_ (.CLK(net183),
    .D(_01054_),
    .Q(\rbzero.tex_b0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21466_ (.CLK(net184),
    .D(_01055_),
    .Q(\rbzero.tex_b0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21467_ (.CLK(net185),
    .D(_01056_),
    .Q(\rbzero.tex_b0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21468_ (.CLK(net186),
    .D(_01057_),
    .Q(\rbzero.tex_b0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21469_ (.CLK(net187),
    .D(_01058_),
    .Q(\rbzero.tex_b0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21470_ (.CLK(net188),
    .D(_01059_),
    .Q(\rbzero.tex_b0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21471_ (.CLK(net189),
    .D(_01060_),
    .Q(\rbzero.tex_b0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21472_ (.CLK(net190),
    .D(_01061_),
    .Q(\rbzero.tex_b0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21473_ (.CLK(net191),
    .D(_01062_),
    .Q(\rbzero.tex_b0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21474_ (.CLK(net192),
    .D(_01063_),
    .Q(\rbzero.tex_b0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21475_ (.CLK(net193),
    .D(_01064_),
    .Q(\rbzero.tex_b0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21476_ (.CLK(net194),
    .D(_01065_),
    .Q(\rbzero.tex_b0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21477_ (.CLK(net195),
    .D(_01066_),
    .Q(\rbzero.tex_b0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21478_ (.CLK(net196),
    .D(_01067_),
    .Q(\rbzero.tex_b0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21479_ (.CLK(net197),
    .D(_01068_),
    .Q(\rbzero.tex_b0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21480_ (.CLK(net198),
    .D(_01069_),
    .Q(\rbzero.tex_b0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21481_ (.CLK(net199),
    .D(_01070_),
    .Q(\rbzero.tex_b0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21482_ (.CLK(net200),
    .D(_01071_),
    .Q(\rbzero.tex_b0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21483_ (.CLK(net201),
    .D(_01072_),
    .Q(\rbzero.tex_b0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21484_ (.CLK(net202),
    .D(_01073_),
    .Q(\rbzero.tex_b0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21485_ (.CLK(net203),
    .D(_01074_),
    .Q(\rbzero.tex_b0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21486_ (.CLK(net204),
    .D(_01075_),
    .Q(\rbzero.tex_b0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21487_ (.CLK(net205),
    .D(_01076_),
    .Q(\rbzero.tex_b0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21488_ (.CLK(net206),
    .D(_01077_),
    .Q(\rbzero.tex_b0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21489_ (.CLK(net207),
    .D(_01078_),
    .Q(\rbzero.tex_b0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21490_ (.CLK(net208),
    .D(_01079_),
    .Q(\rbzero.tex_b0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21491_ (.CLK(net209),
    .D(_01080_),
    .Q(\rbzero.tex_b0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21492_ (.CLK(net210),
    .D(_01081_),
    .Q(\rbzero.tex_b0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21493_ (.CLK(net211),
    .D(_01082_),
    .Q(\rbzero.tex_b0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21494_ (.CLK(net212),
    .D(_01083_),
    .Q(\rbzero.tex_b0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21495_ (.CLK(net213),
    .D(_01084_),
    .Q(\rbzero.tex_b0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21496_ (.CLK(net214),
    .D(_01085_),
    .Q(\rbzero.tex_b0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21497_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01086_),
    .Q(\rbzero.pov.spi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21498_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01087_),
    .Q(\rbzero.pov.spi_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21499_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01088_),
    .Q(\rbzero.pov.spi_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21500_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01089_),
    .Q(\rbzero.pov.spi_buffer[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21501_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01090_),
    .Q(\rbzero.pov.spi_buffer[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21502_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01091_),
    .Q(\rbzero.pov.spi_buffer[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21503_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01092_),
    .Q(\rbzero.pov.spi_buffer[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21504_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01093_),
    .Q(\rbzero.pov.spi_buffer[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21505_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01094_),
    .Q(\rbzero.pov.spi_buffer[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21506_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01095_),
    .Q(\rbzero.pov.spi_buffer[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21507_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01096_),
    .Q(\rbzero.pov.spi_buffer[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21508_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01097_),
    .Q(\rbzero.pov.spi_buffer[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21509_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01098_),
    .Q(\rbzero.pov.spi_buffer[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21510_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01099_),
    .Q(\rbzero.pov.spi_buffer[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21511_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01100_),
    .Q(\rbzero.pov.spi_buffer[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21512_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01101_),
    .Q(\rbzero.pov.spi_buffer[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21513_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01102_),
    .Q(\rbzero.pov.spi_buffer[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21514_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01103_),
    .Q(\rbzero.pov.spi_buffer[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21515_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01104_),
    .Q(\rbzero.pov.spi_buffer[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21516_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01105_),
    .Q(\rbzero.pov.spi_buffer[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21517_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01106_),
    .Q(\rbzero.pov.spi_buffer[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21518_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01107_),
    .Q(\rbzero.pov.spi_buffer[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21519_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01108_),
    .Q(\rbzero.pov.spi_buffer[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21520_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01109_),
    .Q(\rbzero.pov.spi_buffer[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21521_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01110_),
    .Q(\rbzero.pov.spi_buffer[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21522_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01111_),
    .Q(\rbzero.pov.spi_buffer[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21523_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01112_),
    .Q(\rbzero.pov.spi_buffer[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21524_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01113_),
    .Q(\rbzero.pov.spi_buffer[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21525_ (.CLK(clknet_leaf_84_i_clk),
    .D(_01114_),
    .Q(\rbzero.pov.spi_buffer[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21526_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01115_),
    .Q(\rbzero.pov.spi_buffer[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21527_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01116_),
    .Q(\rbzero.pov.spi_buffer[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21528_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01117_),
    .Q(\rbzero.pov.spi_buffer[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21529_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01118_),
    .Q(\rbzero.pov.spi_buffer[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21530_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01119_),
    .Q(\rbzero.pov.spi_buffer[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21531_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01120_),
    .Q(\rbzero.pov.spi_buffer[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21532_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01121_),
    .Q(\rbzero.pov.spi_buffer[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21533_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01122_),
    .Q(\rbzero.pov.spi_buffer[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21534_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01123_),
    .Q(\rbzero.pov.spi_buffer[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21535_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01124_),
    .Q(\rbzero.pov.spi_buffer[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21536_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01125_),
    .Q(\rbzero.pov.spi_buffer[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21537_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01126_),
    .Q(\rbzero.pov.spi_buffer[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21538_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01127_),
    .Q(\rbzero.pov.spi_buffer[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21539_ (.CLK(clknet_leaf_73_i_clk),
    .D(_01128_),
    .Q(\rbzero.pov.spi_buffer[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21540_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01129_),
    .Q(\rbzero.pov.spi_buffer[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21541_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01130_),
    .Q(\rbzero.pov.spi_buffer[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21542_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01131_),
    .Q(\rbzero.pov.spi_buffer[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21543_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01132_),
    .Q(\rbzero.pov.spi_buffer[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21544_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01133_),
    .Q(\rbzero.pov.spi_buffer[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21545_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01134_),
    .Q(\rbzero.pov.spi_buffer[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21546_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01135_),
    .Q(\rbzero.pov.spi_buffer[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21547_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01136_),
    .Q(\rbzero.pov.spi_buffer[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21548_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01137_),
    .Q(\rbzero.pov.spi_buffer[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21549_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01138_),
    .Q(\rbzero.pov.spi_buffer[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21550_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01139_),
    .Q(\rbzero.pov.spi_buffer[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21551_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01140_),
    .Q(\rbzero.pov.spi_buffer[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21552_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01141_),
    .Q(\rbzero.pov.spi_buffer[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21553_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01142_),
    .Q(\rbzero.pov.spi_buffer[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21554_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01143_),
    .Q(\rbzero.pov.spi_buffer[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21555_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01144_),
    .Q(\rbzero.pov.spi_buffer[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21556_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01145_),
    .Q(\rbzero.pov.spi_buffer[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21557_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01146_),
    .Q(\rbzero.pov.spi_buffer[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21558_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01147_),
    .Q(\rbzero.pov.spi_buffer[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21559_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01148_),
    .Q(\rbzero.pov.spi_buffer[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21560_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01149_),
    .Q(\rbzero.pov.spi_buffer[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21561_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01150_),
    .Q(\rbzero.pov.spi_buffer[64] ));
 sky130_fd_sc_hd__dfxtp_1 _21562_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01151_),
    .Q(\rbzero.pov.spi_buffer[65] ));
 sky130_fd_sc_hd__dfxtp_1 _21563_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01152_),
    .Q(\rbzero.pov.spi_buffer[66] ));
 sky130_fd_sc_hd__dfxtp_1 _21564_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01153_),
    .Q(\rbzero.pov.spi_buffer[67] ));
 sky130_fd_sc_hd__dfxtp_1 _21565_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01154_),
    .Q(\rbzero.pov.spi_buffer[68] ));
 sky130_fd_sc_hd__dfxtp_1 _21566_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01155_),
    .Q(\rbzero.pov.spi_buffer[69] ));
 sky130_fd_sc_hd__dfxtp_1 _21567_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01156_),
    .Q(\rbzero.pov.spi_buffer[70] ));
 sky130_fd_sc_hd__dfxtp_1 _21568_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01157_),
    .Q(\rbzero.pov.spi_buffer[71] ));
 sky130_fd_sc_hd__dfxtp_1 _21569_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01158_),
    .Q(\rbzero.pov.spi_buffer[72] ));
 sky130_fd_sc_hd__dfxtp_1 _21570_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01159_),
    .Q(\rbzero.pov.spi_buffer[73] ));
 sky130_fd_sc_hd__dfxtp_1 _21571_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01160_),
    .Q(\rbzero.pov.mosi_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21572_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01161_),
    .Q(\rbzero.pov.mosi ));
 sky130_fd_sc_hd__dfxtp_1 _21573_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01162_),
    .Q(\rbzero.pov.ss_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21574_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01163_),
    .Q(\rbzero.pov.ss_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21575_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01164_),
    .Q(\rbzero.pov.sclk_buffer[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21576_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01165_),
    .Q(\rbzero.pov.sclk_buffer[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21577_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01166_),
    .Q(\rbzero.pov.sclk_buffer[2] ));
 sky130_fd_sc_hd__dfxtp_4 _21578_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01167_),
    .Q(\rbzero.debug_overlay.playerX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21579_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01168_),
    .Q(\rbzero.debug_overlay.playerX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21580_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01169_),
    .Q(\rbzero.debug_overlay.playerX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21581_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01170_),
    .Q(\rbzero.debug_overlay.playerX[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21582_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01171_),
    .Q(\rbzero.debug_overlay.playerX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21583_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01172_),
    .Q(\rbzero.debug_overlay.playerX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21584_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01173_),
    .Q(\rbzero.debug_overlay.playerX[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21585_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01174_),
    .Q(\rbzero.debug_overlay.playerX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21586_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01175_),
    .Q(\rbzero.debug_overlay.playerX[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21587_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01176_),
    .Q(\rbzero.debug_overlay.playerX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21588_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01177_),
    .Q(\rbzero.debug_overlay.playerX[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21589_ (.CLK(clknet_leaf_16_i_clk),
    .D(_01178_),
    .Q(\rbzero.debug_overlay.playerX[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21590_ (.CLK(clknet_leaf_15_i_clk),
    .D(_01179_),
    .Q(\rbzero.debug_overlay.playerX[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21591_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01180_),
    .Q(\rbzero.debug_overlay.playerX[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21592_ (.CLK(clknet_leaf_15_i_clk),
    .D(_01181_),
    .Q(\rbzero.debug_overlay.playerX[5] ));
 sky130_fd_sc_hd__dfxtp_2 _21593_ (.CLK(clknet_leaf_69_i_clk),
    .D(_01182_),
    .Q(\rbzero.debug_overlay.playerY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21594_ (.CLK(clknet_leaf_69_i_clk),
    .D(_01183_),
    .Q(\rbzero.debug_overlay.playerY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21595_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01184_),
    .Q(\rbzero.debug_overlay.playerY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21596_ (.CLK(clknet_leaf_69_i_clk),
    .D(_01185_),
    .Q(\rbzero.debug_overlay.playerY[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21597_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01186_),
    .Q(\rbzero.debug_overlay.playerY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21598_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01187_),
    .Q(\rbzero.debug_overlay.playerY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21599_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01188_),
    .Q(\rbzero.debug_overlay.playerY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21600_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01189_),
    .Q(\rbzero.debug_overlay.playerY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21601_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01190_),
    .Q(\rbzero.debug_overlay.playerY[-1] ));
 sky130_fd_sc_hd__dfxtp_2 _21602_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01191_),
    .Q(\rbzero.debug_overlay.playerY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21603_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01192_),
    .Q(\rbzero.debug_overlay.playerY[1] ));
 sky130_fd_sc_hd__dfxtp_2 _21604_ (.CLK(clknet_leaf_15_i_clk),
    .D(_01193_),
    .Q(\rbzero.debug_overlay.playerY[2] ));
 sky130_fd_sc_hd__dfxtp_2 _21605_ (.CLK(clknet_leaf_13_i_clk),
    .D(_01194_),
    .Q(\rbzero.debug_overlay.playerY[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21606_ (.CLK(clknet_leaf_15_i_clk),
    .D(_01195_),
    .Q(\rbzero.debug_overlay.playerY[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21607_ (.CLK(clknet_leaf_15_i_clk),
    .D(_01196_),
    .Q(\rbzero.debug_overlay.playerY[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21608_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01197_),
    .Q(\rbzero.debug_overlay.facingX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21609_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01198_),
    .Q(\rbzero.debug_overlay.facingX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21610_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01199_),
    .Q(\rbzero.debug_overlay.facingX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21611_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01200_),
    .Q(\rbzero.debug_overlay.facingX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21612_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01201_),
    .Q(\rbzero.debug_overlay.facingX[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21613_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01202_),
    .Q(\rbzero.debug_overlay.facingX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21614_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01203_),
    .Q(\rbzero.debug_overlay.facingX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21615_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01204_),
    .Q(\rbzero.debug_overlay.facingX[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21616_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01205_),
    .Q(\rbzero.debug_overlay.facingX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21617_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01206_),
    .Q(\rbzero.debug_overlay.facingX[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21618_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01207_),
    .Q(\rbzero.debug_overlay.facingX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21619_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01208_),
    .Q(\rbzero.debug_overlay.facingY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _21620_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01209_),
    .Q(\rbzero.debug_overlay.facingY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _21621_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01210_),
    .Q(\rbzero.debug_overlay.facingY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21622_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01211_),
    .Q(\rbzero.debug_overlay.facingY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21623_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01212_),
    .Q(\rbzero.debug_overlay.facingY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21624_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01213_),
    .Q(\rbzero.debug_overlay.facingY[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _21625_ (.CLK(clknet_leaf_87_i_clk),
    .D(_01214_),
    .Q(\rbzero.debug_overlay.facingY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21626_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01215_),
    .Q(\rbzero.debug_overlay.facingY[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _21627_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01216_),
    .Q(\rbzero.debug_overlay.facingY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21628_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01217_),
    .Q(\rbzero.debug_overlay.facingY[0] ));
 sky130_fd_sc_hd__dfxtp_2 _21629_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01218_),
    .Q(\rbzero.debug_overlay.facingY[10] ));
 sky130_fd_sc_hd__dfxtp_4 _21630_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01219_),
    .Q(\rbzero.debug_overlay.vplaneX[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21631_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01220_),
    .Q(\rbzero.debug_overlay.vplaneX[-8] ));
 sky130_fd_sc_hd__dfxtp_4 _21632_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01221_),
    .Q(\rbzero.debug_overlay.vplaneX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21633_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01222_),
    .Q(\rbzero.debug_overlay.vplaneX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _21634_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01223_),
    .Q(\rbzero.debug_overlay.vplaneX[-5] ));
 sky130_fd_sc_hd__dfxtp_4 _21635_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01224_),
    .Q(\rbzero.debug_overlay.vplaneX[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21636_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01225_),
    .Q(\rbzero.debug_overlay.vplaneX[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _21637_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01226_),
    .Q(\rbzero.debug_overlay.vplaneX[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21638_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01227_),
    .Q(\rbzero.debug_overlay.vplaneX[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21639_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01228_),
    .Q(\rbzero.debug_overlay.vplaneX[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21640_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01229_),
    .Q(\rbzero.debug_overlay.vplaneX[10] ));
 sky130_fd_sc_hd__dfxtp_2 _21641_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01230_),
    .Q(\rbzero.debug_overlay.vplaneY[-9] ));
 sky130_fd_sc_hd__dfxtp_2 _21642_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01231_),
    .Q(\rbzero.debug_overlay.vplaneY[-8] ));
 sky130_fd_sc_hd__dfxtp_2 _21643_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01232_),
    .Q(\rbzero.debug_overlay.vplaneY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _21644_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01233_),
    .Q(\rbzero.debug_overlay.vplaneY[-6] ));
 sky130_fd_sc_hd__dfxtp_2 _21645_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01234_),
    .Q(\rbzero.debug_overlay.vplaneY[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _21646_ (.CLK(clknet_leaf_80_i_clk),
    .D(_01235_),
    .Q(\rbzero.debug_overlay.vplaneY[-4] ));
 sky130_fd_sc_hd__dfxtp_2 _21647_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01236_),
    .Q(\rbzero.debug_overlay.vplaneY[-3] ));
 sky130_fd_sc_hd__dfxtp_2 _21648_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01237_),
    .Q(\rbzero.debug_overlay.vplaneY[-2] ));
 sky130_fd_sc_hd__dfxtp_2 _21649_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01238_),
    .Q(\rbzero.debug_overlay.vplaneY[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _21650_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01239_),
    .Q(\rbzero.debug_overlay.vplaneY[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21651_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01240_),
    .Q(\rbzero.debug_overlay.vplaneY[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21652_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01241_),
    .Q(\rbzero.pov.spi_done ));
 sky130_fd_sc_hd__dfxtp_1 _21653_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01242_),
    .Q(\rbzero.vga_sync.vsync ));
 sky130_fd_sc_hd__dfxtp_1 _21654_ (.CLK(clknet_leaf_43_i_clk),
    .D(_01243_),
    .Q(\rbzero.hsync ));
 sky130_fd_sc_hd__dfxtp_2 _21655_ (.CLK(clknet_leaf_44_i_clk),
    .D(_01244_),
    .Q(\gpout0.vpos[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21656_ (.CLK(clknet_leaf_44_i_clk),
    .D(_01245_),
    .Q(\gpout0.vpos[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21657_ (.CLK(clknet_leaf_44_i_clk),
    .D(_01246_),
    .Q(\gpout0.vpos[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21658_ (.CLK(clknet_leaf_17_i_clk),
    .D(_01247_),
    .Q(\gpout0.vpos[3] ));
 sky130_fd_sc_hd__dfxtp_2 _21659_ (.CLK(clknet_leaf_17_i_clk),
    .D(_01248_),
    .Q(\gpout0.vpos[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21660_ (.CLK(clknet_leaf_17_i_clk),
    .D(_01249_),
    .Q(\gpout0.vpos[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21661_ (.CLK(clknet_leaf_19_i_clk),
    .D(_01250_),
    .Q(\gpout0.vpos[6] ));
 sky130_fd_sc_hd__dfxtp_2 _21662_ (.CLK(clknet_leaf_19_i_clk),
    .D(_01251_),
    .Q(\gpout0.vpos[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21663_ (.CLK(clknet_leaf_19_i_clk),
    .D(_01252_),
    .Q(\gpout0.vpos[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21664_ (.CLK(clknet_leaf_19_i_clk),
    .D(_01253_),
    .Q(\gpout0.vpos[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21665_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01254_),
    .Q(\rbzero.spi_registers.new_texadd[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _21666_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01255_),
    .Q(\rbzero.spi_registers.new_texadd[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _21667_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01256_),
    .Q(\rbzero.spi_registers.new_texadd[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _21668_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01257_),
    .Q(\rbzero.spi_registers.new_texadd[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _21669_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01258_),
    .Q(\rbzero.spi_registers.new_texadd[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _21670_ (.CLK(clknet_leaf_31_i_clk),
    .D(_01259_),
    .Q(\rbzero.spi_registers.new_texadd[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _21671_ (.CLK(clknet_leaf_25_i_clk),
    .D(_01260_),
    .Q(\rbzero.spi_registers.new_texadd[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _21672_ (.CLK(clknet_leaf_26_i_clk),
    .D(_01261_),
    .Q(\rbzero.spi_registers.new_texadd[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _21673_ (.CLK(clknet_leaf_7_i_clk),
    .D(_01262_),
    .Q(\rbzero.spi_registers.new_texadd[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _21674_ (.CLK(clknet_leaf_7_i_clk),
    .D(_01263_),
    .Q(\rbzero.spi_registers.new_texadd[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _21675_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01264_),
    .Q(\rbzero.spi_registers.new_texadd[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _21676_ (.CLK(clknet_leaf_0_i_clk),
    .D(_01265_),
    .Q(\rbzero.spi_registers.new_texadd[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _21677_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01266_),
    .Q(\rbzero.spi_registers.new_texadd[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _21678_ (.CLK(clknet_leaf_1_i_clk),
    .D(_01267_),
    .Q(\rbzero.spi_registers.new_texadd[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _21679_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01268_),
    .Q(\rbzero.spi_registers.new_texadd[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _21680_ (.CLK(clknet_leaf_0_i_clk),
    .D(_01269_),
    .Q(\rbzero.spi_registers.new_texadd[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _21681_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01270_),
    .Q(\rbzero.spi_registers.new_texadd[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _21682_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01271_),
    .Q(\rbzero.spi_registers.new_texadd[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _21683_ (.CLK(clknet_leaf_3_i_clk),
    .D(_01272_),
    .Q(\rbzero.spi_registers.new_texadd[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _21684_ (.CLK(clknet_leaf_3_i_clk),
    .D(_01273_),
    .Q(\rbzero.spi_registers.new_texadd[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _21685_ (.CLK(clknet_leaf_3_i_clk),
    .D(_01274_),
    .Q(\rbzero.spi_registers.new_texadd[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _21686_ (.CLK(clknet_leaf_3_i_clk),
    .D(_01275_),
    .Q(\rbzero.spi_registers.new_texadd[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _21687_ (.CLK(clknet_leaf_6_i_clk),
    .D(_01276_),
    .Q(\rbzero.spi_registers.new_texadd[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _21688_ (.CLK(clknet_leaf_6_i_clk),
    .D(_01277_),
    .Q(\rbzero.spi_registers.new_texadd[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _21689_ (.CLK(net215),
    .D(_01278_),
    .Q(\rbzero.tex_b1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21690_ (.CLK(net216),
    .D(_01279_),
    .Q(\rbzero.tex_b1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21691_ (.CLK(net217),
    .D(_01280_),
    .Q(\rbzero.tex_b1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21692_ (.CLK(net218),
    .D(_01281_),
    .Q(\rbzero.tex_b1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21693_ (.CLK(net219),
    .D(_01282_),
    .Q(\rbzero.tex_b1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21694_ (.CLK(net220),
    .D(_01283_),
    .Q(\rbzero.tex_b1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21695_ (.CLK(net221),
    .D(_01284_),
    .Q(\rbzero.tex_b1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21696_ (.CLK(net222),
    .D(_01285_),
    .Q(\rbzero.tex_b1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21697_ (.CLK(net223),
    .D(_01286_),
    .Q(\rbzero.tex_b1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21698_ (.CLK(net224),
    .D(_01287_),
    .Q(\rbzero.tex_b1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21699_ (.CLK(net225),
    .D(_01288_),
    .Q(\rbzero.tex_b1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21700_ (.CLK(net226),
    .D(_01289_),
    .Q(\rbzero.tex_b1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21701_ (.CLK(net227),
    .D(_01290_),
    .Q(\rbzero.tex_b1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21702_ (.CLK(net228),
    .D(_01291_),
    .Q(\rbzero.tex_b1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21703_ (.CLK(net229),
    .D(_01292_),
    .Q(\rbzero.tex_b1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21704_ (.CLK(net230),
    .D(_01293_),
    .Q(\rbzero.tex_b1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21705_ (.CLK(net231),
    .D(_01294_),
    .Q(\rbzero.tex_b1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21706_ (.CLK(net232),
    .D(_01295_),
    .Q(\rbzero.tex_b1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21707_ (.CLK(net233),
    .D(_01296_),
    .Q(\rbzero.tex_b1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21708_ (.CLK(net234),
    .D(_01297_),
    .Q(\rbzero.tex_b1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21709_ (.CLK(net235),
    .D(_01298_),
    .Q(\rbzero.tex_b1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21710_ (.CLK(net236),
    .D(_01299_),
    .Q(\rbzero.tex_b1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21711_ (.CLK(net237),
    .D(_01300_),
    .Q(\rbzero.tex_b1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21712_ (.CLK(net238),
    .D(_01301_),
    .Q(\rbzero.tex_b1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21713_ (.CLK(net239),
    .D(_01302_),
    .Q(\rbzero.tex_b1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21714_ (.CLK(net240),
    .D(_01303_),
    .Q(\rbzero.tex_b1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21715_ (.CLK(net241),
    .D(_01304_),
    .Q(\rbzero.tex_b1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21716_ (.CLK(net242),
    .D(_01305_),
    .Q(\rbzero.tex_b1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21717_ (.CLK(net243),
    .D(_01306_),
    .Q(\rbzero.tex_b1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21718_ (.CLK(net244),
    .D(_01307_),
    .Q(\rbzero.tex_b1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21719_ (.CLK(net245),
    .D(_01308_),
    .Q(\rbzero.tex_b1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21720_ (.CLK(net246),
    .D(_01309_),
    .Q(\rbzero.tex_b1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21721_ (.CLK(net247),
    .D(_01310_),
    .Q(\rbzero.tex_b1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21722_ (.CLK(net248),
    .D(_01311_),
    .Q(\rbzero.tex_b1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21723_ (.CLK(net249),
    .D(_01312_),
    .Q(\rbzero.tex_b1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21724_ (.CLK(net250),
    .D(_01313_),
    .Q(\rbzero.tex_b1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21725_ (.CLK(net251),
    .D(_01314_),
    .Q(\rbzero.tex_b1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21726_ (.CLK(net252),
    .D(_01315_),
    .Q(\rbzero.tex_b1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21727_ (.CLK(net253),
    .D(_01316_),
    .Q(\rbzero.tex_b1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21728_ (.CLK(net254),
    .D(_01317_),
    .Q(\rbzero.tex_b1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21729_ (.CLK(net255),
    .D(_01318_),
    .Q(\rbzero.tex_b1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21730_ (.CLK(net256),
    .D(_01319_),
    .Q(\rbzero.tex_b1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21731_ (.CLK(net257),
    .D(_01320_),
    .Q(\rbzero.tex_b1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21732_ (.CLK(net258),
    .D(_01321_),
    .Q(\rbzero.tex_b1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21733_ (.CLK(net259),
    .D(_01322_),
    .Q(\rbzero.tex_b1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21734_ (.CLK(net260),
    .D(_01323_),
    .Q(\rbzero.tex_b1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21735_ (.CLK(net261),
    .D(_01324_),
    .Q(\rbzero.tex_b1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21736_ (.CLK(net262),
    .D(_01325_),
    .Q(\rbzero.tex_b1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21737_ (.CLK(net263),
    .D(_01326_),
    .Q(\rbzero.tex_b1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21738_ (.CLK(net264),
    .D(_01327_),
    .Q(\rbzero.tex_b1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21739_ (.CLK(net265),
    .D(_01328_),
    .Q(\rbzero.tex_b1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21740_ (.CLK(net266),
    .D(_01329_),
    .Q(\rbzero.tex_b1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21741_ (.CLK(net267),
    .D(_01330_),
    .Q(\rbzero.tex_b1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21742_ (.CLK(net268),
    .D(_01331_),
    .Q(\rbzero.tex_b1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21743_ (.CLK(net269),
    .D(_01332_),
    .Q(\rbzero.tex_b1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21744_ (.CLK(net270),
    .D(_01333_),
    .Q(\rbzero.tex_b1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21745_ (.CLK(net271),
    .D(_01334_),
    .Q(\rbzero.tex_b1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21746_ (.CLK(net272),
    .D(_01335_),
    .Q(\rbzero.tex_b1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21747_ (.CLK(net273),
    .D(_01336_),
    .Q(\rbzero.tex_b1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21748_ (.CLK(net274),
    .D(_01337_),
    .Q(\rbzero.tex_b1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21749_ (.CLK(net275),
    .D(_01338_),
    .Q(\rbzero.tex_b1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21750_ (.CLK(net276),
    .D(_01339_),
    .Q(\rbzero.tex_b1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21751_ (.CLK(net277),
    .D(_01340_),
    .Q(\rbzero.tex_b1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21752_ (.CLK(net278),
    .D(_01341_),
    .Q(\rbzero.tex_b1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21753_ (.CLK(net279),
    .D(_01342_),
    .Q(\rbzero.tex_g0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21754_ (.CLK(net280),
    .D(_01343_),
    .Q(\rbzero.tex_g0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21755_ (.CLK(net281),
    .D(_01344_),
    .Q(\rbzero.tex_g0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21756_ (.CLK(net282),
    .D(_01345_),
    .Q(\rbzero.tex_g0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21757_ (.CLK(net283),
    .D(_01346_),
    .Q(\rbzero.tex_g0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21758_ (.CLK(net284),
    .D(_01347_),
    .Q(\rbzero.tex_g0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21759_ (.CLK(net285),
    .D(_01348_),
    .Q(\rbzero.tex_g0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21760_ (.CLK(net286),
    .D(_01349_),
    .Q(\rbzero.tex_g0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21761_ (.CLK(net287),
    .D(_01350_),
    .Q(\rbzero.tex_g0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21762_ (.CLK(net288),
    .D(_01351_),
    .Q(\rbzero.tex_g0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21763_ (.CLK(net289),
    .D(_01352_),
    .Q(\rbzero.tex_g0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21764_ (.CLK(net290),
    .D(_01353_),
    .Q(\rbzero.tex_g0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21765_ (.CLK(net291),
    .D(_01354_),
    .Q(\rbzero.tex_g0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21766_ (.CLK(net292),
    .D(_01355_),
    .Q(\rbzero.tex_g0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21767_ (.CLK(net293),
    .D(_01356_),
    .Q(\rbzero.tex_g0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21768_ (.CLK(net294),
    .D(_01357_),
    .Q(\rbzero.tex_g0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21769_ (.CLK(net295),
    .D(_01358_),
    .Q(\rbzero.tex_g0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21770_ (.CLK(net296),
    .D(_01359_),
    .Q(\rbzero.tex_g0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21771_ (.CLK(net297),
    .D(_01360_),
    .Q(\rbzero.tex_g0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21772_ (.CLK(net298),
    .D(_01361_),
    .Q(\rbzero.tex_g0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21773_ (.CLK(net299),
    .D(_01362_),
    .Q(\rbzero.tex_g0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21774_ (.CLK(net300),
    .D(_01363_),
    .Q(\rbzero.tex_g0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21775_ (.CLK(net301),
    .D(_01364_),
    .Q(\rbzero.tex_g0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21776_ (.CLK(net302),
    .D(_01365_),
    .Q(\rbzero.tex_g0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21777_ (.CLK(net303),
    .D(_01366_),
    .Q(\rbzero.tex_g0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21778_ (.CLK(net304),
    .D(_01367_),
    .Q(\rbzero.tex_g0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21779_ (.CLK(net305),
    .D(_01368_),
    .Q(\rbzero.tex_g0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21780_ (.CLK(net306),
    .D(_01369_),
    .Q(\rbzero.tex_g0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21781_ (.CLK(net307),
    .D(_01370_),
    .Q(\rbzero.tex_g0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21782_ (.CLK(net308),
    .D(_01371_),
    .Q(\rbzero.tex_g0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21783_ (.CLK(net309),
    .D(_01372_),
    .Q(\rbzero.tex_g0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21784_ (.CLK(net310),
    .D(_01373_),
    .Q(\rbzero.tex_g0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21785_ (.CLK(net311),
    .D(_01374_),
    .Q(\rbzero.tex_g0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21786_ (.CLK(net312),
    .D(_01375_),
    .Q(\rbzero.tex_g0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21787_ (.CLK(net313),
    .D(_01376_),
    .Q(\rbzero.tex_g0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21788_ (.CLK(net314),
    .D(_01377_),
    .Q(\rbzero.tex_g0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21789_ (.CLK(net315),
    .D(_01378_),
    .Q(\rbzero.tex_g0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21790_ (.CLK(net316),
    .D(_01379_),
    .Q(\rbzero.tex_g0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21791_ (.CLK(net317),
    .D(_01380_),
    .Q(\rbzero.tex_g0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21792_ (.CLK(net318),
    .D(_01381_),
    .Q(\rbzero.tex_g0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21793_ (.CLK(net319),
    .D(_01382_),
    .Q(\rbzero.tex_g0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21794_ (.CLK(net320),
    .D(_01383_),
    .Q(\rbzero.tex_g0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21795_ (.CLK(net321),
    .D(_01384_),
    .Q(\rbzero.tex_g0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21796_ (.CLK(net322),
    .D(_01385_),
    .Q(\rbzero.tex_g0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21797_ (.CLK(net323),
    .D(_01386_),
    .Q(\rbzero.tex_g0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21798_ (.CLK(net324),
    .D(_01387_),
    .Q(\rbzero.tex_g0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21799_ (.CLK(net325),
    .D(_01388_),
    .Q(\rbzero.tex_g0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21800_ (.CLK(net326),
    .D(_01389_),
    .Q(\rbzero.tex_g0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21801_ (.CLK(net327),
    .D(_01390_),
    .Q(\rbzero.tex_g0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21802_ (.CLK(net328),
    .D(_01391_),
    .Q(\rbzero.tex_g0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21803_ (.CLK(net329),
    .D(_01392_),
    .Q(\rbzero.tex_g0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21804_ (.CLK(net330),
    .D(_01393_),
    .Q(\rbzero.tex_g0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21805_ (.CLK(net331),
    .D(_01394_),
    .Q(\rbzero.tex_g0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21806_ (.CLK(net332),
    .D(_01395_),
    .Q(\rbzero.tex_g0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21807_ (.CLK(net333),
    .D(_01396_),
    .Q(\rbzero.tex_g0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21808_ (.CLK(net334),
    .D(_01397_),
    .Q(\rbzero.tex_g0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21809_ (.CLK(net335),
    .D(_01398_),
    .Q(\rbzero.tex_g0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21810_ (.CLK(net336),
    .D(_01399_),
    .Q(\rbzero.tex_g0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21811_ (.CLK(net337),
    .D(_01400_),
    .Q(\rbzero.tex_g0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21812_ (.CLK(net338),
    .D(_01401_),
    .Q(\rbzero.tex_g0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21813_ (.CLK(net339),
    .D(_01402_),
    .Q(\rbzero.tex_g0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21814_ (.CLK(net340),
    .D(_01403_),
    .Q(\rbzero.tex_g0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21815_ (.CLK(net341),
    .D(_01404_),
    .Q(\rbzero.tex_g0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21816_ (.CLK(net342),
    .D(_01405_),
    .Q(\rbzero.tex_g0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21817_ (.CLK(net343),
    .D(_01406_),
    .Q(\rbzero.tex_g1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21818_ (.CLK(net344),
    .D(_01407_),
    .Q(\rbzero.tex_g1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21819_ (.CLK(net345),
    .D(_01408_),
    .Q(\rbzero.tex_g1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21820_ (.CLK(net346),
    .D(_01409_),
    .Q(\rbzero.tex_g1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21821_ (.CLK(net347),
    .D(_01410_),
    .Q(\rbzero.tex_g1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21822_ (.CLK(net348),
    .D(_01411_),
    .Q(\rbzero.tex_g1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21823_ (.CLK(net349),
    .D(_01412_),
    .Q(\rbzero.tex_g1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21824_ (.CLK(net350),
    .D(_01413_),
    .Q(\rbzero.tex_g1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21825_ (.CLK(net351),
    .D(_01414_),
    .Q(\rbzero.tex_g1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21826_ (.CLK(net352),
    .D(_01415_),
    .Q(\rbzero.tex_g1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21827_ (.CLK(net353),
    .D(_01416_),
    .Q(\rbzero.tex_g1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21828_ (.CLK(net354),
    .D(_01417_),
    .Q(\rbzero.tex_g1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21829_ (.CLK(net355),
    .D(_01418_),
    .Q(\rbzero.tex_g1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21830_ (.CLK(net356),
    .D(_01419_),
    .Q(\rbzero.tex_g1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21831_ (.CLK(net357),
    .D(_01420_),
    .Q(\rbzero.tex_g1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21832_ (.CLK(net358),
    .D(_01421_),
    .Q(\rbzero.tex_g1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21833_ (.CLK(net359),
    .D(_01422_),
    .Q(\rbzero.tex_g1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21834_ (.CLK(net360),
    .D(_01423_),
    .Q(\rbzero.tex_g1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21835_ (.CLK(net361),
    .D(_01424_),
    .Q(\rbzero.tex_g1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21836_ (.CLK(net362),
    .D(_01425_),
    .Q(\rbzero.tex_g1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21837_ (.CLK(net363),
    .D(_01426_),
    .Q(\rbzero.tex_g1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21838_ (.CLK(net364),
    .D(_01427_),
    .Q(\rbzero.tex_g1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21839_ (.CLK(net365),
    .D(_01428_),
    .Q(\rbzero.tex_g1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21840_ (.CLK(net366),
    .D(_01429_),
    .Q(\rbzero.tex_g1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21841_ (.CLK(net367),
    .D(_01430_),
    .Q(\rbzero.tex_g1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21842_ (.CLK(net368),
    .D(_01431_),
    .Q(\rbzero.tex_g1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21843_ (.CLK(net369),
    .D(_01432_),
    .Q(\rbzero.tex_g1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21844_ (.CLK(net370),
    .D(_01433_),
    .Q(\rbzero.tex_g1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21845_ (.CLK(net371),
    .D(_01434_),
    .Q(\rbzero.tex_g1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21846_ (.CLK(net372),
    .D(_01435_),
    .Q(\rbzero.tex_g1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21847_ (.CLK(net373),
    .D(_01436_),
    .Q(\rbzero.tex_g1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21848_ (.CLK(net374),
    .D(_01437_),
    .Q(\rbzero.tex_g1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21849_ (.CLK(net375),
    .D(_01438_),
    .Q(\rbzero.tex_g1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21850_ (.CLK(net376),
    .D(_01439_),
    .Q(\rbzero.tex_g1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21851_ (.CLK(net377),
    .D(_01440_),
    .Q(\rbzero.tex_g1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21852_ (.CLK(net378),
    .D(_01441_),
    .Q(\rbzero.tex_g1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21853_ (.CLK(net379),
    .D(_01442_),
    .Q(\rbzero.tex_g1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21854_ (.CLK(net380),
    .D(_01443_),
    .Q(\rbzero.tex_g1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21855_ (.CLK(net381),
    .D(_01444_),
    .Q(\rbzero.tex_g1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21856_ (.CLK(net382),
    .D(_01445_),
    .Q(\rbzero.tex_g1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21857_ (.CLK(net383),
    .D(_01446_),
    .Q(\rbzero.tex_g1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21858_ (.CLK(net384),
    .D(_01447_),
    .Q(\rbzero.tex_g1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21859_ (.CLK(net385),
    .D(_01448_),
    .Q(\rbzero.tex_g1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21860_ (.CLK(net386),
    .D(_01449_),
    .Q(\rbzero.tex_g1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21861_ (.CLK(net387),
    .D(_01450_),
    .Q(\rbzero.tex_g1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21862_ (.CLK(net388),
    .D(_01451_),
    .Q(\rbzero.tex_g1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21863_ (.CLK(net389),
    .D(_01452_),
    .Q(\rbzero.tex_g1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21864_ (.CLK(net390),
    .D(_01453_),
    .Q(\rbzero.tex_g1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21865_ (.CLK(net391),
    .D(_01454_),
    .Q(\rbzero.tex_g1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21866_ (.CLK(net392),
    .D(_01455_),
    .Q(\rbzero.tex_g1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21867_ (.CLK(net393),
    .D(_01456_),
    .Q(\rbzero.tex_g1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21868_ (.CLK(net394),
    .D(_01457_),
    .Q(\rbzero.tex_g1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21869_ (.CLK(net395),
    .D(_01458_),
    .Q(\rbzero.tex_g1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21870_ (.CLK(net396),
    .D(_01459_),
    .Q(\rbzero.tex_g1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21871_ (.CLK(net397),
    .D(_01460_),
    .Q(\rbzero.tex_g1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21872_ (.CLK(net398),
    .D(_01461_),
    .Q(\rbzero.tex_g1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21873_ (.CLK(net399),
    .D(_01462_),
    .Q(\rbzero.tex_g1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21874_ (.CLK(net400),
    .D(_01463_),
    .Q(\rbzero.tex_g1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21875_ (.CLK(net401),
    .D(_01464_),
    .Q(\rbzero.tex_g1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21876_ (.CLK(net402),
    .D(_01465_),
    .Q(\rbzero.tex_g1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21877_ (.CLK(net403),
    .D(_01466_),
    .Q(\rbzero.tex_g1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21878_ (.CLK(net404),
    .D(_01467_),
    .Q(\rbzero.tex_g1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21879_ (.CLK(net405),
    .D(_01468_),
    .Q(\rbzero.tex_g1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21880_ (.CLK(net406),
    .D(_01469_),
    .Q(\rbzero.tex_g1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21881_ (.CLK(net407),
    .D(_01470_),
    .Q(\rbzero.tex_r0[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21882_ (.CLK(net408),
    .D(_01471_),
    .Q(\rbzero.tex_r0[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21883_ (.CLK(net409),
    .D(_01472_),
    .Q(\rbzero.tex_r0[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21884_ (.CLK(net410),
    .D(_01473_),
    .Q(\rbzero.tex_r0[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21885_ (.CLK(net411),
    .D(_01474_),
    .Q(\rbzero.tex_r0[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21886_ (.CLK(net412),
    .D(_01475_),
    .Q(\rbzero.tex_r0[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21887_ (.CLK(net413),
    .D(_01476_),
    .Q(\rbzero.tex_r0[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21888_ (.CLK(net414),
    .D(_01477_),
    .Q(\rbzero.tex_r0[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21889_ (.CLK(net415),
    .D(_01478_),
    .Q(\rbzero.tex_r0[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21890_ (.CLK(net416),
    .D(_01479_),
    .Q(\rbzero.tex_r0[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21891_ (.CLK(net417),
    .D(_01480_),
    .Q(\rbzero.tex_r0[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21892_ (.CLK(net418),
    .D(_01481_),
    .Q(\rbzero.tex_r0[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21893_ (.CLK(net419),
    .D(_01482_),
    .Q(\rbzero.tex_r0[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21894_ (.CLK(net420),
    .D(_01483_),
    .Q(\rbzero.tex_r0[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21895_ (.CLK(net421),
    .D(_01484_),
    .Q(\rbzero.tex_r0[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21896_ (.CLK(net422),
    .D(_01485_),
    .Q(\rbzero.tex_r0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21897_ (.CLK(net423),
    .D(_01486_),
    .Q(\rbzero.tex_r0[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21898_ (.CLK(net424),
    .D(_01487_),
    .Q(\rbzero.tex_r0[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21899_ (.CLK(net425),
    .D(_01488_),
    .Q(\rbzero.tex_r0[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21900_ (.CLK(net426),
    .D(_01489_),
    .Q(\rbzero.tex_r0[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21901_ (.CLK(net427),
    .D(_01490_),
    .Q(\rbzero.tex_r0[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21902_ (.CLK(net428),
    .D(_01491_),
    .Q(\rbzero.tex_r0[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21903_ (.CLK(net429),
    .D(_01492_),
    .Q(\rbzero.tex_r0[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21904_ (.CLK(net430),
    .D(_01493_),
    .Q(\rbzero.tex_r0[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21905_ (.CLK(net431),
    .D(_01494_),
    .Q(\rbzero.tex_r0[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21906_ (.CLK(net432),
    .D(_01495_),
    .Q(\rbzero.tex_r0[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21907_ (.CLK(net433),
    .D(_01496_),
    .Q(\rbzero.tex_r0[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21908_ (.CLK(net434),
    .D(_01497_),
    .Q(\rbzero.tex_r0[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21909_ (.CLK(net435),
    .D(_01498_),
    .Q(\rbzero.tex_r0[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21910_ (.CLK(net436),
    .D(_01499_),
    .Q(\rbzero.tex_r0[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21911_ (.CLK(net437),
    .D(_01500_),
    .Q(\rbzero.tex_r0[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21912_ (.CLK(net438),
    .D(_01501_),
    .Q(\rbzero.tex_r0[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21913_ (.CLK(net439),
    .D(_01502_),
    .Q(\rbzero.tex_r0[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21914_ (.CLK(net440),
    .D(_01503_),
    .Q(\rbzero.tex_r0[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21915_ (.CLK(net441),
    .D(_01504_),
    .Q(\rbzero.tex_r0[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21916_ (.CLK(net442),
    .D(_01505_),
    .Q(\rbzero.tex_r0[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21917_ (.CLK(net443),
    .D(_01506_),
    .Q(\rbzero.tex_r0[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21918_ (.CLK(net444),
    .D(_01507_),
    .Q(\rbzero.tex_r0[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21919_ (.CLK(net445),
    .D(_01508_),
    .Q(\rbzero.tex_r0[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21920_ (.CLK(net446),
    .D(_01509_),
    .Q(\rbzero.tex_r0[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21921_ (.CLK(net447),
    .D(_01510_),
    .Q(\rbzero.tex_r0[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21922_ (.CLK(net448),
    .D(_01511_),
    .Q(\rbzero.tex_r0[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21923_ (.CLK(net449),
    .D(_01512_),
    .Q(\rbzero.tex_r0[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21924_ (.CLK(net450),
    .D(_01513_),
    .Q(\rbzero.tex_r0[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21925_ (.CLK(net451),
    .D(_01514_),
    .Q(\rbzero.tex_r0[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21926_ (.CLK(net452),
    .D(_01515_),
    .Q(\rbzero.tex_r0[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21927_ (.CLK(net453),
    .D(_01516_),
    .Q(\rbzero.tex_r0[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21928_ (.CLK(net454),
    .D(_01517_),
    .Q(\rbzero.tex_r0[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21929_ (.CLK(net455),
    .D(_01518_),
    .Q(\rbzero.tex_r0[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21930_ (.CLK(net456),
    .D(_01519_),
    .Q(\rbzero.tex_r0[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21931_ (.CLK(net457),
    .D(_01520_),
    .Q(\rbzero.tex_r0[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21932_ (.CLK(net458),
    .D(_01521_),
    .Q(\rbzero.tex_r0[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21933_ (.CLK(net459),
    .D(_01522_),
    .Q(\rbzero.tex_r0[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21934_ (.CLK(net460),
    .D(_01523_),
    .Q(\rbzero.tex_r0[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21935_ (.CLK(net461),
    .D(_01524_),
    .Q(\rbzero.tex_r0[54] ));
 sky130_fd_sc_hd__dfxtp_1 _21936_ (.CLK(net462),
    .D(_01525_),
    .Q(\rbzero.tex_r0[55] ));
 sky130_fd_sc_hd__dfxtp_1 _21937_ (.CLK(net463),
    .D(_01526_),
    .Q(\rbzero.tex_r0[56] ));
 sky130_fd_sc_hd__dfxtp_1 _21938_ (.CLK(net464),
    .D(_01527_),
    .Q(\rbzero.tex_r0[57] ));
 sky130_fd_sc_hd__dfxtp_1 _21939_ (.CLK(net465),
    .D(_01528_),
    .Q(\rbzero.tex_r0[58] ));
 sky130_fd_sc_hd__dfxtp_1 _21940_ (.CLK(net466),
    .D(_01529_),
    .Q(\rbzero.tex_r0[59] ));
 sky130_fd_sc_hd__dfxtp_1 _21941_ (.CLK(net467),
    .D(_01530_),
    .Q(\rbzero.tex_r0[60] ));
 sky130_fd_sc_hd__dfxtp_1 _21942_ (.CLK(net468),
    .D(_01531_),
    .Q(\rbzero.tex_r0[61] ));
 sky130_fd_sc_hd__dfxtp_1 _21943_ (.CLK(net469),
    .D(_01532_),
    .Q(\rbzero.tex_r0[62] ));
 sky130_fd_sc_hd__dfxtp_1 _21944_ (.CLK(net470),
    .D(_01533_),
    .Q(\rbzero.tex_r0[63] ));
 sky130_fd_sc_hd__dfxtp_1 _21945_ (.CLK(net471),
    .D(_01534_),
    .Q(\rbzero.tex_r1[0] ));
 sky130_fd_sc_hd__dfxtp_1 _21946_ (.CLK(net472),
    .D(_01535_),
    .Q(\rbzero.tex_r1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _21947_ (.CLK(net473),
    .D(_01536_),
    .Q(\rbzero.tex_r1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _21948_ (.CLK(net474),
    .D(_01537_),
    .Q(\rbzero.tex_r1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _21949_ (.CLK(net475),
    .D(_01538_),
    .Q(\rbzero.tex_r1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _21950_ (.CLK(net476),
    .D(_01539_),
    .Q(\rbzero.tex_r1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _21951_ (.CLK(net477),
    .D(_01540_),
    .Q(\rbzero.tex_r1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _21952_ (.CLK(net478),
    .D(_01541_),
    .Q(\rbzero.tex_r1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _21953_ (.CLK(net479),
    .D(_01542_),
    .Q(\rbzero.tex_r1[8] ));
 sky130_fd_sc_hd__dfxtp_1 _21954_ (.CLK(net480),
    .D(_01543_),
    .Q(\rbzero.tex_r1[9] ));
 sky130_fd_sc_hd__dfxtp_1 _21955_ (.CLK(net481),
    .D(_01544_),
    .Q(\rbzero.tex_r1[10] ));
 sky130_fd_sc_hd__dfxtp_1 _21956_ (.CLK(net482),
    .D(_01545_),
    .Q(\rbzero.tex_r1[11] ));
 sky130_fd_sc_hd__dfxtp_1 _21957_ (.CLK(net483),
    .D(_01546_),
    .Q(\rbzero.tex_r1[12] ));
 sky130_fd_sc_hd__dfxtp_1 _21958_ (.CLK(net484),
    .D(_01547_),
    .Q(\rbzero.tex_r1[13] ));
 sky130_fd_sc_hd__dfxtp_1 _21959_ (.CLK(net485),
    .D(_01548_),
    .Q(\rbzero.tex_r1[14] ));
 sky130_fd_sc_hd__dfxtp_1 _21960_ (.CLK(net486),
    .D(_01549_),
    .Q(\rbzero.tex_r1[15] ));
 sky130_fd_sc_hd__dfxtp_1 _21961_ (.CLK(net487),
    .D(_01550_),
    .Q(\rbzero.tex_r1[16] ));
 sky130_fd_sc_hd__dfxtp_1 _21962_ (.CLK(net488),
    .D(_01551_),
    .Q(\rbzero.tex_r1[17] ));
 sky130_fd_sc_hd__dfxtp_1 _21963_ (.CLK(net489),
    .D(_01552_),
    .Q(\rbzero.tex_r1[18] ));
 sky130_fd_sc_hd__dfxtp_1 _21964_ (.CLK(net490),
    .D(_01553_),
    .Q(\rbzero.tex_r1[19] ));
 sky130_fd_sc_hd__dfxtp_1 _21965_ (.CLK(net491),
    .D(_01554_),
    .Q(\rbzero.tex_r1[20] ));
 sky130_fd_sc_hd__dfxtp_1 _21966_ (.CLK(net492),
    .D(_01555_),
    .Q(\rbzero.tex_r1[21] ));
 sky130_fd_sc_hd__dfxtp_1 _21967_ (.CLK(net493),
    .D(_01556_),
    .Q(\rbzero.tex_r1[22] ));
 sky130_fd_sc_hd__dfxtp_1 _21968_ (.CLK(net494),
    .D(_01557_),
    .Q(\rbzero.tex_r1[23] ));
 sky130_fd_sc_hd__dfxtp_1 _21969_ (.CLK(net495),
    .D(_01558_),
    .Q(\rbzero.tex_r1[24] ));
 sky130_fd_sc_hd__dfxtp_1 _21970_ (.CLK(net496),
    .D(_01559_),
    .Q(\rbzero.tex_r1[25] ));
 sky130_fd_sc_hd__dfxtp_1 _21971_ (.CLK(net497),
    .D(_01560_),
    .Q(\rbzero.tex_r1[26] ));
 sky130_fd_sc_hd__dfxtp_1 _21972_ (.CLK(net498),
    .D(_01561_),
    .Q(\rbzero.tex_r1[27] ));
 sky130_fd_sc_hd__dfxtp_1 _21973_ (.CLK(net499),
    .D(_01562_),
    .Q(\rbzero.tex_r1[28] ));
 sky130_fd_sc_hd__dfxtp_1 _21974_ (.CLK(net500),
    .D(_01563_),
    .Q(\rbzero.tex_r1[29] ));
 sky130_fd_sc_hd__dfxtp_1 _21975_ (.CLK(net501),
    .D(_01564_),
    .Q(\rbzero.tex_r1[30] ));
 sky130_fd_sc_hd__dfxtp_1 _21976_ (.CLK(net502),
    .D(_01565_),
    .Q(\rbzero.tex_r1[31] ));
 sky130_fd_sc_hd__dfxtp_1 _21977_ (.CLK(net503),
    .D(_01566_),
    .Q(\rbzero.tex_r1[32] ));
 sky130_fd_sc_hd__dfxtp_1 _21978_ (.CLK(net504),
    .D(_01567_),
    .Q(\rbzero.tex_r1[33] ));
 sky130_fd_sc_hd__dfxtp_1 _21979_ (.CLK(net505),
    .D(_01568_),
    .Q(\rbzero.tex_r1[34] ));
 sky130_fd_sc_hd__dfxtp_1 _21980_ (.CLK(net506),
    .D(_01569_),
    .Q(\rbzero.tex_r1[35] ));
 sky130_fd_sc_hd__dfxtp_1 _21981_ (.CLK(net507),
    .D(_01570_),
    .Q(\rbzero.tex_r1[36] ));
 sky130_fd_sc_hd__dfxtp_1 _21982_ (.CLK(net508),
    .D(_01571_),
    .Q(\rbzero.tex_r1[37] ));
 sky130_fd_sc_hd__dfxtp_1 _21983_ (.CLK(net509),
    .D(_01572_),
    .Q(\rbzero.tex_r1[38] ));
 sky130_fd_sc_hd__dfxtp_1 _21984_ (.CLK(net510),
    .D(_01573_),
    .Q(\rbzero.tex_r1[39] ));
 sky130_fd_sc_hd__dfxtp_1 _21985_ (.CLK(net131),
    .D(_01574_),
    .Q(\rbzero.tex_r1[40] ));
 sky130_fd_sc_hd__dfxtp_1 _21986_ (.CLK(net132),
    .D(_01575_),
    .Q(\rbzero.tex_r1[41] ));
 sky130_fd_sc_hd__dfxtp_1 _21987_ (.CLK(net133),
    .D(_01576_),
    .Q(\rbzero.tex_r1[42] ));
 sky130_fd_sc_hd__dfxtp_1 _21988_ (.CLK(net134),
    .D(_01577_),
    .Q(\rbzero.tex_r1[43] ));
 sky130_fd_sc_hd__dfxtp_1 _21989_ (.CLK(net135),
    .D(_01578_),
    .Q(\rbzero.tex_r1[44] ));
 sky130_fd_sc_hd__dfxtp_1 _21990_ (.CLK(net136),
    .D(_01579_),
    .Q(\rbzero.tex_r1[45] ));
 sky130_fd_sc_hd__dfxtp_1 _21991_ (.CLK(net137),
    .D(_01580_),
    .Q(\rbzero.tex_r1[46] ));
 sky130_fd_sc_hd__dfxtp_1 _21992_ (.CLK(net138),
    .D(_01581_),
    .Q(\rbzero.tex_r1[47] ));
 sky130_fd_sc_hd__dfxtp_1 _21993_ (.CLK(net139),
    .D(_01582_),
    .Q(\rbzero.tex_r1[48] ));
 sky130_fd_sc_hd__dfxtp_1 _21994_ (.CLK(net140),
    .D(_01583_),
    .Q(\rbzero.tex_r1[49] ));
 sky130_fd_sc_hd__dfxtp_1 _21995_ (.CLK(net141),
    .D(_01584_),
    .Q(\rbzero.tex_r1[50] ));
 sky130_fd_sc_hd__dfxtp_1 _21996_ (.CLK(net142),
    .D(_01585_),
    .Q(\rbzero.tex_r1[51] ));
 sky130_fd_sc_hd__dfxtp_1 _21997_ (.CLK(net143),
    .D(_01586_),
    .Q(\rbzero.tex_r1[52] ));
 sky130_fd_sc_hd__dfxtp_1 _21998_ (.CLK(net144),
    .D(_01587_),
    .Q(\rbzero.tex_r1[53] ));
 sky130_fd_sc_hd__dfxtp_1 _21999_ (.CLK(net145),
    .D(_01588_),
    .Q(\rbzero.tex_r1[54] ));
 sky130_fd_sc_hd__dfxtp_1 _22000_ (.CLK(net146),
    .D(_01589_),
    .Q(\rbzero.tex_r1[55] ));
 sky130_fd_sc_hd__dfxtp_1 _22001_ (.CLK(net147),
    .D(_01590_),
    .Q(\rbzero.tex_r1[56] ));
 sky130_fd_sc_hd__dfxtp_1 _22002_ (.CLK(net148),
    .D(_01591_),
    .Q(\rbzero.tex_r1[57] ));
 sky130_fd_sc_hd__dfxtp_1 _22003_ (.CLK(net149),
    .D(_01592_),
    .Q(\rbzero.tex_r1[58] ));
 sky130_fd_sc_hd__dfxtp_1 _22004_ (.CLK(net150),
    .D(_01593_),
    .Q(\rbzero.tex_r1[59] ));
 sky130_fd_sc_hd__dfxtp_1 _22005_ (.CLK(net127),
    .D(_01594_),
    .Q(\rbzero.tex_r1[60] ));
 sky130_fd_sc_hd__dfxtp_1 _22006_ (.CLK(net128),
    .D(_01595_),
    .Q(\rbzero.tex_r1[61] ));
 sky130_fd_sc_hd__dfxtp_1 _22007_ (.CLK(net129),
    .D(_01596_),
    .Q(\rbzero.tex_r1[62] ));
 sky130_fd_sc_hd__dfxtp_1 _22008_ (.CLK(net130),
    .D(_01597_),
    .Q(\rbzero.tex_r1[63] ));
 sky130_fd_sc_hd__dfxtp_1 _22009_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01598_),
    .Q(\gpout5.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22010_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01599_),
    .Q(\gpout5.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22011_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01600_),
    .Q(\rbzero.texV[-11] ));
 sky130_fd_sc_hd__dfxtp_1 _22012_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01601_),
    .Q(\rbzero.texV[-10] ));
 sky130_fd_sc_hd__dfxtp_1 _22013_ (.CLK(clknet_leaf_68_i_clk),
    .D(_01602_),
    .Q(\rbzero.texV[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22014_ (.CLK(clknet_leaf_69_i_clk),
    .D(_01603_),
    .Q(\rbzero.texV[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22015_ (.CLK(clknet_leaf_48_i_clk),
    .D(_01604_),
    .Q(\rbzero.texV[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22016_ (.CLK(clknet_leaf_69_i_clk),
    .D(_01605_),
    .Q(\rbzero.texV[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22017_ (.CLK(clknet_leaf_48_i_clk),
    .D(_01606_),
    .Q(\rbzero.texV[-5] ));
 sky130_fd_sc_hd__dfxtp_1 _22018_ (.CLK(clknet_leaf_48_i_clk),
    .D(_01607_),
    .Q(\rbzero.texV[-4] ));
 sky130_fd_sc_hd__dfxtp_1 _22019_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01608_),
    .Q(\rbzero.texV[-3] ));
 sky130_fd_sc_hd__dfxtp_1 _22020_ (.CLK(clknet_leaf_49_i_clk),
    .D(_01609_),
    .Q(\rbzero.texV[-2] ));
 sky130_fd_sc_hd__dfxtp_1 _22021_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01610_),
    .Q(\rbzero.texV[-1] ));
 sky130_fd_sc_hd__dfxtp_1 _22022_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01611_),
    .Q(\rbzero.texV[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22023_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01612_),
    .Q(\rbzero.texV[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22024_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01613_),
    .Q(\rbzero.texV[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22025_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01614_),
    .Q(\rbzero.texV[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22026_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01615_),
    .Q(\rbzero.texV[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22027_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01616_),
    .Q(\rbzero.texV[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22028_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01617_),
    .Q(\rbzero.texV[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22029_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01618_),
    .Q(\rbzero.texV[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22030_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01619_),
    .Q(\rbzero.texV[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22031_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01620_),
    .Q(\rbzero.texV[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22032_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01621_),
    .Q(\rbzero.texV[10] ));
 sky130_fd_sc_hd__dfxtp_4 _22033_ (.CLK(clknet_leaf_67_i_clk),
    .D(_01622_),
    .Q(\rbzero.trace_state[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22034_ (.CLK(clknet_leaf_67_i_clk),
    .D(_01623_),
    .Q(\rbzero.trace_state[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22035_ (.CLK(clknet_leaf_68_i_clk),
    .D(_01624_),
    .Q(\rbzero.trace_state[2] ));
 sky130_fd_sc_hd__dfxtp_4 _22036_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01625_),
    .Q(\rbzero.trace_state[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22037_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01626_),
    .Q(\reg_gpout[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22038_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01627_),
    .Q(\reg_gpout[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22039_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01628_),
    .Q(\reg_gpout[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22040_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01629_),
    .Q(\reg_gpout[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22041_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01630_),
    .Q(\reg_gpout[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22042_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01631_),
    .Q(\reg_gpout[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22043_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01632_),
    .Q(reg_hsync));
 sky130_fd_sc_hd__dfxtp_1 _22044_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01633_),
    .Q(reg_vsync));
 sky130_fd_sc_hd__dfxtp_1 _22045_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01634_),
    .Q(\rbzero.traced_texVinit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22046_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01635_),
    .Q(\rbzero.traced_texVinit[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22047_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01636_),
    .Q(\rbzero.traced_texVinit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _22048_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01637_),
    .Q(\rbzero.traced_texVinit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _22049_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01638_),
    .Q(\rbzero.traced_texVinit[4] ));
 sky130_fd_sc_hd__dfxtp_1 _22050_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01639_),
    .Q(\rbzero.traced_texVinit[5] ));
 sky130_fd_sc_hd__dfxtp_1 _22051_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01640_),
    .Q(\rbzero.traced_texVinit[6] ));
 sky130_fd_sc_hd__dfxtp_1 _22052_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01641_),
    .Q(\rbzero.traced_texVinit[7] ));
 sky130_fd_sc_hd__dfxtp_1 _22053_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01642_),
    .Q(\rbzero.traced_texVinit[8] ));
 sky130_fd_sc_hd__dfxtp_1 _22054_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01643_),
    .Q(\rbzero.traced_texVinit[9] ));
 sky130_fd_sc_hd__dfxtp_1 _22055_ (.CLK(clknet_leaf_54_i_clk),
    .D(_01644_),
    .Q(\rbzero.traced_texVinit[10] ));
 sky130_fd_sc_hd__dfxtp_1 _22056_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01645_),
    .Q(\gpout0.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22057_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01646_),
    .Q(\gpout0.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22058_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01647_),
    .Q(\rbzero.wall_tracer.rayAddendX[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22059_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01648_),
    .Q(\rbzero.wall_tracer.rayAddendX[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22060_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01649_),
    .Q(\rbzero.wall_tracer.rayAddendX[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22061_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01650_),
    .Q(\rbzero.wall_tracer.rayAddendX[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22062_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01651_),
    .Q(\rbzero.wall_tracer.rayAddendY[-9] ));
 sky130_fd_sc_hd__dfxtp_1 _22063_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01652_),
    .Q(\rbzero.wall_tracer.rayAddendY[-8] ));
 sky130_fd_sc_hd__dfxtp_1 _22064_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01653_),
    .Q(\rbzero.wall_tracer.rayAddendY[-7] ));
 sky130_fd_sc_hd__dfxtp_1 _22065_ (.CLK(clknet_leaf_79_i_clk),
    .D(_01654_),
    .Q(\rbzero.wall_tracer.rayAddendY[-6] ));
 sky130_fd_sc_hd__dfxtp_1 _22066_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01655_),
    .Q(\gpout1.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22067_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01656_),
    .Q(\gpout1.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22068_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01657_),
    .Q(\gpout2.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22069_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01658_),
    .Q(\gpout2.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22070_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01659_),
    .Q(\gpout3.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22071_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01660_),
    .Q(\gpout3.clk_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _22072_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01661_),
    .Q(\gpout4.clk_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _22073_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01662_),
    .Q(\gpout4.clk_div[1] ));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_110 (.HI(net110));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_111 (.HI(net111));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_112 (.HI(net112));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_113 (.HI(net113));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_114 (.HI(net114));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_115 (.HI(net115));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_116 (.HI(net116));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_117 (.HI(net117));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_118 (.HI(net118));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_119 (.HI(net119));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_120 (.HI(net120));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_121 (.HI(net121));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_122 (.HI(net122));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_123 (.HI(net123));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_124 (.HI(net124));
 sky130_fd_sc_hd__inv_2 _11444__1 (.A(clknet_1_1__leaf__04634_),
    .Y(net125));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_76 (.LO(net76));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_77 (.LO(net77));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_78 (.LO(net78));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_79 (.LO(net79));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_80 (.LO(net80));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_81 (.LO(net81));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_82 (.LO(net82));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_83 (.LO(net83));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_84 (.LO(net84));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_85 (.LO(net85));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_86 (.LO(net86));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_87 (.LO(net87));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_88 (.LO(net88));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_89 (.LO(net89));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_90 (.LO(net90));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_91 (.LO(net91));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_92 (.LO(net92));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_93 (.LO(net93));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_94 (.LO(net94));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_95 (.LO(net95));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_96 (.LO(net96));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_99 (.LO(net99));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_100 (.LO(net100));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_101 (.LO(net101));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_102 (.LO(net102));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_103 (.LO(net103));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_104 (.LO(net104));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_105 (.LO(net105));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_106 (.LO(net106));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_107 (.LO(net107));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_108 (.LO(net108));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_109 (.HI(net109));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(i_debug_map_overlay),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(i_debug_trace_overlay),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(i_debug_vec_overlay),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input4 (.A(i_gpout0_sel[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_6 input5 (.A(i_gpout0_sel[1]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(i_gpout0_sel[2]),
    .X(net6));
 sky130_fd_sc_hd__buf_6 input7 (.A(i_gpout0_sel[3]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(i_gpout0_sel[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(i_gpout0_sel[5]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input10 (.A(i_gpout1_sel[0]),
    .X(net10));
 sky130_fd_sc_hd__buf_6 input11 (.A(i_gpout1_sel[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_8 input12 (.A(i_gpout1_sel[2]),
    .X(net12));
 sky130_fd_sc_hd__buf_6 input13 (.A(i_gpout1_sel[3]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_8 input14 (.A(i_gpout1_sel[4]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(i_gpout1_sel[5]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input16 (.A(i_gpout2_sel[0]),
    .X(net16));
 sky130_fd_sc_hd__buf_6 input17 (.A(i_gpout2_sel[1]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(i_gpout2_sel[2]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input19 (.A(i_gpout2_sel[3]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input20 (.A(i_gpout2_sel[4]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input21 (.A(i_gpout2_sel[5]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input22 (.A(i_gpout3_sel[0]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_8 input23 (.A(i_gpout3_sel[1]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(i_gpout3_sel[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_8 input25 (.A(i_gpout3_sel[3]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(i_gpout3_sel[4]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(i_gpout3_sel[5]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(i_gpout4_sel[0]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(i_gpout4_sel[1]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 input30 (.A(i_gpout4_sel[2]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(i_gpout4_sel[3]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(i_gpout4_sel[4]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(i_gpout4_sel[5]),
    .X(net33));
 sky130_fd_sc_hd__buf_6 input34 (.A(i_gpout5_sel[0]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(i_gpout5_sel[1]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(i_gpout5_sel[2]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(i_gpout5_sel[3]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(i_gpout5_sel[4]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(i_gpout5_sel[5]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_16 input40 (.A(i_mode[0]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_16 input41 (.A(i_mode[1]),
    .X(net41));
 sky130_fd_sc_hd__buf_4 input42 (.A(i_mode[2]),
    .X(net42));
 sky130_fd_sc_hd__buf_8 input43 (.A(i_reg_csb),
    .X(net43));
 sky130_fd_sc_hd__buf_8 input44 (.A(i_reg_mosi),
    .X(net44));
 sky130_fd_sc_hd__buf_6 input45 (.A(i_reg_outs_enb),
    .X(net45));
 sky130_fd_sc_hd__buf_6 input46 (.A(i_reg_sclk),
    .X(net46));
 sky130_fd_sc_hd__buf_4 input47 (.A(i_reset_lock_a),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_8 input48 (.A(i_reset_lock_b),
    .X(net48));
 sky130_fd_sc_hd__buf_6 input49 (.A(i_tex_in[0]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 input50 (.A(i_tex_in[1]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 input51 (.A(i_tex_in[2]),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(i_tex_in[3]),
    .X(net52));
 sky130_fd_sc_hd__buf_6 input53 (.A(i_vec_csb),
    .X(net53));
 sky130_fd_sc_hd__buf_4 input54 (.A(i_vec_mosi),
    .X(net54));
 sky130_fd_sc_hd__buf_6 input55 (.A(i_vec_sclk),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(o_gpout[0]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(o_gpout[1]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(o_gpout[2]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(o_gpout[3]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(o_gpout[4]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(o_gpout[5]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(o_hsync));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(o_reset));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(o_rgb[14]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(o_rgb[15]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(o_rgb[22]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(o_rgb[23]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(o_rgb[6]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(o_rgb[7]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(o_tex_csb));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(o_tex_oeb0));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(o_tex_out0));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net125),
    .X(o_tex_sclk));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(o_vsync));
 sky130_fd_sc_hd__conb_1 top_ew_algofoogle_75 (.LO(net75));
 sky130_fd_sc_hd__inv_2 net99_2 (.A(clknet_1_0__leaf__04634_),
    .Y(net126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_opt_2_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_opt_3_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_opt_4_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_51_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_52_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_53_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_54_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_55_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_56_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_57_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_58_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_59_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_60_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_61_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_62_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_63_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_64_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_65_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_66_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_leaf_67_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_leaf_68_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_69_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_70_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_71_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_72_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_73_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_74_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_76_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_77_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_78_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_79_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_80_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_81_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_82_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_83_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_84_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_85_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_leaf_86_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_87_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_88_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_89_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_leaf_90_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_91_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_92_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_93_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_94_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_95_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_96_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_leaf_97_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_i_clk (.A(clknet_opt_1_0_i_clk),
    .X(clknet_leaf_98_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_99_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_leaf_100_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_opt_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_2_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_opt_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_3_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_opt_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_4_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_opt_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05820_ (.A(_05820_),
    .X(clknet_0__05820_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05820_ (.A(clknet_0__05820_),
    .X(clknet_1_0__leaf__05820_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05820_ (.A(clknet_0__05820_),
    .X(clknet_1_1__leaf__05820_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05700_ (.A(_05700_),
    .X(clknet_0__05700_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05700_ (.A(clknet_0__05700_),
    .X(clknet_1_0__leaf__05700_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05700_ (.A(clknet_0__05700_),
    .X(clknet_1_1__leaf__05700_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04634_ (.A(_04634_),
    .X(clknet_0__04634_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04634_ (.A(clknet_0__04634_),
    .X(clknet_1_0__leaf__04634_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04634_ (.A(clknet_0__04634_),
    .X(clknet_1_1__leaf__04634_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05993_ (.A(_05993_),
    .X(clknet_0__05993_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05993_ (.A(clknet_0__05993_),
    .X(clknet_1_0__leaf__05993_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05993_ (.A(clknet_0__05993_),
    .X(clknet_1_1__leaf__05993_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03808_ (.A(_03808_),
    .X(clknet_0__03808_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03808_ (.A(clknet_0__03808_),
    .X(clknet_1_0__leaf__03808_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03808_ (.A(clknet_0__03808_),
    .X(clknet_1_1__leaf__03808_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03807_ (.A(_03807_),
    .X(clknet_0__03807_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03807_ (.A(clknet_0__03807_),
    .X(clknet_1_0__leaf__03807_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03807_ (.A(clknet_0__03807_),
    .X(clknet_1_1__leaf__03807_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03796_ (.A(_03796_),
    .X(clknet_0__03796_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03796_ (.A(clknet_0__03796_),
    .X(clknet_1_0__leaf__03796_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03796_ (.A(clknet_0__03796_),
    .X(clknet_1_1__leaf__03796_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03806_ (.A(_03806_),
    .X(clknet_0__03806_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03806_ (.A(clknet_0__03806_),
    .X(clknet_1_0__leaf__03806_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03806_ (.A(clknet_0__03806_),
    .X(clknet_1_1__leaf__03806_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03805_ (.A(_03805_),
    .X(clknet_0__03805_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03805_ (.A(clknet_0__03805_),
    .X(clknet_1_0__leaf__03805_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03805_ (.A(clknet_0__03805_),
    .X(clknet_1_1__leaf__03805_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03804_ (.A(_03804_),
    .X(clknet_0__03804_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03804_ (.A(clknet_0__03804_),
    .X(clknet_1_0__leaf__03804_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03804_ (.A(clknet_0__03804_),
    .X(clknet_1_1__leaf__03804_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03803_ (.A(_03803_),
    .X(clknet_0__03803_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03803_ (.A(clknet_0__03803_),
    .X(clknet_1_0__leaf__03803_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03803_ (.A(clknet_0__03803_),
    .X(clknet_1_1__leaf__03803_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03802_ (.A(_03802_),
    .X(clknet_0__03802_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03802_ (.A(clknet_0__03802_),
    .X(clknet_1_0__leaf__03802_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03802_ (.A(clknet_0__03802_),
    .X(clknet_1_1__leaf__03802_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03801_ (.A(_03801_),
    .X(clknet_0__03801_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03801_ (.A(clknet_0__03801_),
    .X(clknet_1_0__leaf__03801_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03801_ (.A(clknet_0__03801_),
    .X(clknet_1_1__leaf__03801_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03800_ (.A(_03800_),
    .X(clknet_0__03800_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03800_ (.A(clknet_0__03800_),
    .X(clknet_1_0__leaf__03800_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03800_ (.A(clknet_0__03800_),
    .X(clknet_1_1__leaf__03800_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03799_ (.A(_03799_),
    .X(clknet_0__03799_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03799_ (.A(clknet_0__03799_),
    .X(clknet_1_0__leaf__03799_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03799_ (.A(clknet_0__03799_),
    .X(clknet_1_1__leaf__03799_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03798_ (.A(_03798_),
    .X(clknet_0__03798_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03798_ (.A(clknet_0__03798_),
    .X(clknet_1_0__leaf__03798_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03798_ (.A(clknet_0__03798_),
    .X(clknet_1_1__leaf__03798_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03797_ (.A(_03797_),
    .X(clknet_0__03797_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03797_ (.A(clknet_0__03797_),
    .X(clknet_1_0__leaf__03797_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03797_ (.A(clknet_0__03797_),
    .X(clknet_1_1__leaf__03797_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03785_ (.A(_03785_),
    .X(clknet_0__03785_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03785_ (.A(clknet_0__03785_),
    .X(clknet_1_0__leaf__03785_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03785_ (.A(clknet_0__03785_),
    .X(clknet_1_1__leaf__03785_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03795_ (.A(_03795_),
    .X(clknet_0__03795_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03795_ (.A(clknet_0__03795_),
    .X(clknet_1_0__leaf__03795_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03795_ (.A(clknet_0__03795_),
    .X(clknet_1_1__leaf__03795_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03794_ (.A(_03794_),
    .X(clknet_0__03794_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03794_ (.A(clknet_0__03794_),
    .X(clknet_1_0__leaf__03794_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03794_ (.A(clknet_0__03794_),
    .X(clknet_1_1__leaf__03794_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03793_ (.A(_03793_),
    .X(clknet_0__03793_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03793_ (.A(clknet_0__03793_),
    .X(clknet_1_0__leaf__03793_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03793_ (.A(clknet_0__03793_),
    .X(clknet_1_1__leaf__03793_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03792_ (.A(_03792_),
    .X(clknet_0__03792_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03792_ (.A(clknet_0__03792_),
    .X(clknet_1_0__leaf__03792_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03792_ (.A(clknet_0__03792_),
    .X(clknet_1_1__leaf__03792_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03791_ (.A(_03791_),
    .X(clknet_0__03791_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03791_ (.A(clknet_0__03791_),
    .X(clknet_1_0__leaf__03791_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03791_ (.A(clknet_0__03791_),
    .X(clknet_1_1__leaf__03791_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03790_ (.A(_03790_),
    .X(clknet_0__03790_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03790_ (.A(clknet_0__03790_),
    .X(clknet_1_0__leaf__03790_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03790_ (.A(clknet_0__03790_),
    .X(clknet_1_1__leaf__03790_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03789_ (.A(_03789_),
    .X(clknet_0__03789_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03789_ (.A(clknet_0__03789_),
    .X(clknet_1_0__leaf__03789_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03789_ (.A(clknet_0__03789_),
    .X(clknet_1_1__leaf__03789_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03788_ (.A(_03788_),
    .X(clknet_0__03788_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03788_ (.A(clknet_0__03788_),
    .X(clknet_1_0__leaf__03788_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03788_ (.A(clknet_0__03788_),
    .X(clknet_1_1__leaf__03788_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03787_ (.A(_03787_),
    .X(clknet_0__03787_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03787_ (.A(clknet_0__03787_),
    .X(clknet_1_0__leaf__03787_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03787_ (.A(clknet_0__03787_),
    .X(clknet_1_1__leaf__03787_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03786_ (.A(_03786_),
    .X(clknet_0__03786_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03786_ (.A(clknet_0__03786_),
    .X(clknet_1_0__leaf__03786_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03786_ (.A(clknet_0__03786_),
    .X(clknet_1_1__leaf__03786_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03464_ (.A(_03464_),
    .X(clknet_0__03464_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03464_ (.A(clknet_0__03464_),
    .X(clknet_1_0__leaf__03464_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03464_ (.A(clknet_0__03464_),
    .X(clknet_1_1__leaf__03464_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03784_ (.A(_03784_),
    .X(clknet_0__03784_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03784_ (.A(clknet_0__03784_),
    .X(clknet_1_0__leaf__03784_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03784_ (.A(clknet_0__03784_),
    .X(clknet_1_1__leaf__03784_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03783_ (.A(_03783_),
    .X(clknet_0__03783_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03783_ (.A(clknet_0__03783_),
    .X(clknet_1_0__leaf__03783_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03783_ (.A(clknet_0__03783_),
    .X(clknet_1_1__leaf__03783_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03782_ (.A(_03782_),
    .X(clknet_0__03782_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03782_ (.A(clknet_0__03782_),
    .X(clknet_1_0__leaf__03782_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03782_ (.A(clknet_0__03782_),
    .X(clknet_1_1__leaf__03782_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03781_ (.A(_03781_),
    .X(clknet_0__03781_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03781_ (.A(clknet_0__03781_),
    .X(clknet_1_0__leaf__03781_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03781_ (.A(clknet_0__03781_),
    .X(clknet_1_1__leaf__03781_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03780_ (.A(_03780_),
    .X(clknet_0__03780_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03780_ (.A(clknet_0__03780_),
    .X(clknet_1_0__leaf__03780_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03780_ (.A(clknet_0__03780_),
    .X(clknet_1_1__leaf__03780_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03779_ (.A(_03779_),
    .X(clknet_0__03779_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03779_ (.A(clknet_0__03779_),
    .X(clknet_1_0__leaf__03779_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03779_ (.A(clknet_0__03779_),
    .X(clknet_1_1__leaf__03779_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03778_ (.A(_03778_),
    .X(clknet_0__03778_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03778_ (.A(clknet_0__03778_),
    .X(clknet_1_0__leaf__03778_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03778_ (.A(clknet_0__03778_),
    .X(clknet_1_1__leaf__03778_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03777_ (.A(_03777_),
    .X(clknet_0__03777_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03777_ (.A(clknet_0__03777_),
    .X(clknet_1_0__leaf__03777_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03777_ (.A(clknet_0__03777_),
    .X(clknet_1_1__leaf__03777_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03776_ (.A(_03776_),
    .X(clknet_0__03776_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03776_ (.A(clknet_0__03776_),
    .X(clknet_1_0__leaf__03776_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03776_ (.A(clknet_0__03776_),
    .X(clknet_1_1__leaf__03776_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03465_ (.A(_03465_),
    .X(clknet_0__03465_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03465_ (.A(clknet_0__03465_),
    .X(clknet_1_0__leaf__03465_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03465_ (.A(clknet_0__03465_),
    .X(clknet_1_1__leaf__03465_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03457_ (.A(_03457_),
    .X(clknet_0__03457_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03457_ (.A(clknet_0__03457_),
    .X(clknet_1_0__leaf__03457_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03457_ (.A(clknet_0__03457_),
    .X(clknet_1_1__leaf__03457_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03463_ (.A(_03463_),
    .X(clknet_0__03463_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03463_ (.A(clknet_0__03463_),
    .X(clknet_1_0__leaf__03463_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03463_ (.A(clknet_0__03463_),
    .X(clknet_1_1__leaf__03463_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03462_ (.A(_03462_),
    .X(clknet_0__03462_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03462_ (.A(clknet_0__03462_),
    .X(clknet_1_0__leaf__03462_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03462_ (.A(clknet_0__03462_),
    .X(clknet_1_1__leaf__03462_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03461_ (.A(_03461_),
    .X(clknet_0__03461_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03461_ (.A(clknet_0__03461_),
    .X(clknet_1_0__leaf__03461_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03461_ (.A(clknet_0__03461_),
    .X(clknet_1_1__leaf__03461_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03460_ (.A(_03460_),
    .X(clknet_0__03460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03460_ (.A(clknet_0__03460_),
    .X(clknet_1_0__leaf__03460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03460_ (.A(clknet_0__03460_),
    .X(clknet_1_1__leaf__03460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03459_ (.A(_03459_),
    .X(clknet_0__03459_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03459_ (.A(clknet_0__03459_),
    .X(clknet_1_0__leaf__03459_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03459_ (.A(clknet_0__03459_),
    .X(clknet_1_1__leaf__03459_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__03458_ (.A(_03458_),
    .X(clknet_0__03458_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__03458_ (.A(clknet_0__03458_),
    .X(clknet_1_0__leaf__03458_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__03458_ (.A(clknet_0__03458_),
    .X(clknet_1_1__leaf__03458_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05938_ (.A(_05938_),
    .X(clknet_0__05938_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05938_ (.A(clknet_0__05938_),
    .X(clknet_1_0__leaf__05938_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05938_ (.A(clknet_0__05938_),
    .X(clknet_1_1__leaf__05938_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05879_ (.A(_05879_),
    .X(clknet_0__05879_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05879_ (.A(clknet_0__05879_),
    .X(clknet_1_0__leaf__05879_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05879_ (.A(clknet_0__05879_),
    .X(clknet_1_1__leaf__05879_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__05761_ (.A(_05761_),
    .X(clknet_0__05761_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__05761_ (.A(clknet_0__05761_),
    .X(clknet_1_0__leaf__05761_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__05761_ (.A(clknet_0__05761_),
    .X(clknet_1_1__leaf__05761_));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\rbzero.tex_r1[40] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\rbzero.pov.spi_buffer[6] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\rbzero.pov.ready_buffer[43] ),
    .X(net512));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_04429_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_04429_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_04464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_04464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_05064_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_05126_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_05552_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_07935_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_07971_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_08039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_08124_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_08136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_08136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_08136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_08148_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_09747_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_09747_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\rbzero.spi_registers.vshift[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\rbzero.spi_registers.vshift[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\rbzero.tex_r0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\rbzero.trace_state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\rbzero.trace_state[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\rbzero.wall_tracer.visualWallDist[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\rbzero.wall_tracer.visualWallDist[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\rbzero.wall_tracer.visualWallDist[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_05299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_05821_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_07996_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_03110_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net70));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1066 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1120 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1235 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1167 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1094 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1235 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1242 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1078 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1248 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1126 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1176 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1194 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1232 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1222 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1180 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1223 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1143 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1067 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1227 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1240 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1150 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1058 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1066 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1206 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1064 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1070 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1150 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1248 ();
 assign o_rgb[0] = net75;
 assign o_rgb[10] = net83;
 assign o_rgb[11] = net84;
 assign o_rgb[12] = net85;
 assign o_rgb[13] = net86;
 assign o_rgb[16] = net87;
 assign o_rgb[17] = net88;
 assign o_rgb[18] = net89;
 assign o_rgb[19] = net90;
 assign o_rgb[1] = net76;
 assign o_rgb[20] = net91;
 assign o_rgb[21] = net92;
 assign o_rgb[2] = net77;
 assign o_rgb[3] = net78;
 assign o_rgb[4] = net79;
 assign o_rgb[5] = net80;
 assign o_rgb[8] = net81;
 assign o_rgb[9] = net82;
 assign ones[0] = net109;
 assign ones[10] = net119;
 assign ones[11] = net120;
 assign ones[12] = net121;
 assign ones[13] = net122;
 assign ones[14] = net123;
 assign ones[15] = net124;
 assign ones[1] = net110;
 assign ones[2] = net111;
 assign ones[3] = net112;
 assign ones[4] = net113;
 assign ones[5] = net114;
 assign ones[6] = net115;
 assign ones[7] = net116;
 assign ones[8] = net117;
 assign ones[9] = net118;
 assign zeros[0] = net93;
 assign zeros[10] = net103;
 assign zeros[11] = net104;
 assign zeros[12] = net105;
 assign zeros[13] = net106;
 assign zeros[14] = net107;
 assign zeros[15] = net108;
 assign zeros[1] = net94;
 assign zeros[2] = net95;
 assign zeros[3] = net96;
 assign zeros[4] = net97;
 assign zeros[5] = net98;
 assign zeros[6] = net99;
 assign zeros[7] = net100;
 assign zeros[8] = net101;
 assign zeros[9] = net102;
endmodule


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_io_control
  CLASS BLOCK ;
  FOREIGN analog_io_control ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 240.000 ;
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 20.440 80.000 21.040 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 59.880 80.000 60.480 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 99.320 80.000 99.920 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 138.760 80.000 139.360 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 178.200 80.000 178.800 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 76.000 217.640 80.000 218.240 ;
    END
  END io_oeb[5]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 13.285 10.640 14.885 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 30.420 10.640 32.020 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.555 10.640 49.155 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.690 10.640 66.290 228.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.850 10.640 23.450 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.985 10.640 40.585 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.120 10.640 57.720 228.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.255 10.640 74.855 228.720 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 224.345 74.250 227.175 ;
        RECT 5.330 218.905 74.250 221.735 ;
        RECT 5.330 213.465 74.250 216.295 ;
        RECT 5.330 208.025 74.250 210.855 ;
        RECT 5.330 202.585 74.250 205.415 ;
        RECT 5.330 197.145 74.250 199.975 ;
        RECT 5.330 191.705 74.250 194.535 ;
        RECT 5.330 186.265 74.250 189.095 ;
        RECT 5.330 180.825 74.250 183.655 ;
        RECT 5.330 175.385 74.250 178.215 ;
        RECT 5.330 169.945 74.250 172.775 ;
        RECT 5.330 164.505 74.250 167.335 ;
        RECT 5.330 159.065 74.250 161.895 ;
        RECT 5.330 153.625 74.250 156.455 ;
        RECT 5.330 148.185 74.250 151.015 ;
        RECT 5.330 142.745 74.250 145.575 ;
        RECT 5.330 137.305 74.250 140.135 ;
        RECT 5.330 131.865 74.250 134.695 ;
        RECT 5.330 126.425 74.250 129.255 ;
        RECT 5.330 120.985 74.250 123.815 ;
        RECT 5.330 115.545 74.250 118.375 ;
        RECT 5.330 110.105 74.250 112.935 ;
        RECT 5.330 104.665 74.250 107.495 ;
        RECT 5.330 99.225 74.250 102.055 ;
        RECT 5.330 93.785 74.250 96.615 ;
        RECT 5.330 88.345 74.250 91.175 ;
        RECT 5.330 82.905 74.250 85.735 ;
        RECT 5.330 77.465 74.250 80.295 ;
        RECT 5.330 72.025 74.250 74.855 ;
        RECT 5.330 66.585 74.250 69.415 ;
        RECT 5.330 61.145 74.250 63.975 ;
        RECT 5.330 55.705 74.250 58.535 ;
        RECT 5.330 50.265 74.250 53.095 ;
        RECT 5.330 44.825 74.250 47.655 ;
        RECT 5.330 39.385 74.250 42.215 ;
        RECT 5.330 33.945 74.250 36.775 ;
        RECT 5.330 28.505 74.250 31.335 ;
        RECT 5.330 23.065 74.250 25.895 ;
        RECT 5.330 17.625 74.250 20.455 ;
        RECT 5.330 12.185 74.250 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 74.060 228.565 ;
      LAYER met1 ;
        RECT 5.520 10.640 74.855 228.720 ;
      LAYER met2 ;
        RECT 13.315 10.695 74.825 228.665 ;
      LAYER met3 ;
        RECT 13.295 218.640 76.050 228.645 ;
        RECT 13.295 217.240 75.600 218.640 ;
        RECT 13.295 179.200 76.050 217.240 ;
        RECT 13.295 177.800 75.600 179.200 ;
        RECT 13.295 139.760 76.050 177.800 ;
        RECT 13.295 138.360 75.600 139.760 ;
        RECT 13.295 100.320 76.050 138.360 ;
        RECT 13.295 98.920 75.600 100.320 ;
        RECT 13.295 60.880 76.050 98.920 ;
        RECT 13.295 59.480 75.600 60.880 ;
        RECT 13.295 21.440 76.050 59.480 ;
        RECT 13.295 20.040 75.600 21.440 ;
        RECT 13.295 10.715 76.050 20.040 ;
  END
END analog_io_control
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1698657151
<< nwell >>
rect 1066 44869 14850 45435
rect 1066 43781 14850 44347
rect 1066 42693 14850 43259
rect 1066 41605 14850 42171
rect 1066 40517 14850 41083
rect 1066 39429 14850 39995
rect 1066 38341 14850 38907
rect 1066 37253 14850 37819
rect 1066 36165 14850 36731
rect 1066 35077 14850 35643
rect 1066 33989 14850 34555
rect 1066 32901 14850 33467
rect 1066 31813 14850 32379
rect 1066 30725 14850 31291
rect 1066 29637 14850 30203
rect 1066 28549 14850 29115
rect 1066 27461 14850 28027
rect 1066 26373 14850 26939
rect 1066 25285 14850 25851
rect 1066 24197 14850 24763
rect 1066 23109 14850 23675
rect 1066 22021 14850 22587
rect 1066 20933 14850 21499
rect 1066 19845 14850 20411
rect 1066 18757 14850 19323
rect 1066 17669 14850 18235
rect 1066 16581 14850 17147
rect 1066 15493 14850 16059
rect 1066 14405 14850 14971
rect 1066 13317 14850 13883
rect 1066 12229 14850 12795
rect 1066 11141 14850 11707
rect 1066 10053 14850 10619
rect 1066 8965 14850 9531
rect 1066 7877 14850 8443
rect 1066 6789 14850 7355
rect 1066 5701 14850 6267
rect 1066 4613 14850 5179
rect 1066 3525 14850 4091
rect 1066 2437 14850 3003
<< obsli1 >>
rect 1104 2159 14812 45713
<< obsm1 >>
rect 1104 2128 14971 45744
<< obsm2 >>
rect 2663 2139 14965 45733
<< metal3 >>
rect 15200 43528 16000 43648
rect 15200 35640 16000 35760
rect 15200 27752 16000 27872
rect 15200 19864 16000 19984
rect 15200 11976 16000 12096
rect 15200 4088 16000 4208
<< obsm3 >>
rect 2659 43728 15210 45729
rect 2659 43448 15120 43728
rect 2659 35840 15210 43448
rect 2659 35560 15120 35840
rect 2659 27952 15210 35560
rect 2659 27672 15120 27952
rect 2659 20064 15210 27672
rect 2659 19784 15120 20064
rect 2659 12176 15210 19784
rect 2659 11896 15120 12176
rect 2659 4288 15210 11896
rect 2659 4008 15120 4288
rect 2659 2143 15210 4008
<< metal4 >>
rect 2657 2128 2977 45744
rect 4370 2128 4690 45744
rect 6084 2128 6404 45744
rect 7797 2128 8117 45744
rect 9511 2128 9831 45744
rect 11224 2128 11544 45744
rect 12938 2128 13258 45744
rect 14651 2128 14971 45744
<< labels >>
rlabel metal3 s 15200 4088 16000 4208 6 io_oeb[0]
port 1 nsew signal output
rlabel metal3 s 15200 11976 16000 12096 6 io_oeb[1]
port 2 nsew signal output
rlabel metal3 s 15200 19864 16000 19984 6 io_oeb[2]
port 3 nsew signal output
rlabel metal3 s 15200 27752 16000 27872 6 io_oeb[3]
port 4 nsew signal output
rlabel metal3 s 15200 35640 16000 35760 6 io_oeb[4]
port 5 nsew signal output
rlabel metal3 s 15200 43528 16000 43648 6 io_oeb[5]
port 6 nsew signal output
rlabel metal4 s 2657 2128 2977 45744 6 vccd1
port 7 nsew power bidirectional
rlabel metal4 s 6084 2128 6404 45744 6 vccd1
port 7 nsew power bidirectional
rlabel metal4 s 9511 2128 9831 45744 6 vccd1
port 7 nsew power bidirectional
rlabel metal4 s 12938 2128 13258 45744 6 vccd1
port 7 nsew power bidirectional
rlabel metal4 s 4370 2128 4690 45744 6 vssd1
port 8 nsew ground bidirectional
rlabel metal4 s 7797 2128 8117 45744 6 vssd1
port 8 nsew ground bidirectional
rlabel metal4 s 11224 2128 11544 45744 6 vssd1
port 8 nsew ground bidirectional
rlabel metal4 s 14651 2128 14971 45744 6 vssd1
port 8 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 48000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 481330
string GDS_FILE /home/zwierzak/projects/caravel_user_project/openlane/analog_io_control/runs/23_10_30_10_06/results/signoff/analog_io_control.magic.gds
string GDS_START 23768
<< end >>

